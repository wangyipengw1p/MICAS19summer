`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 11/07/2018 11:41:44 AM
// Design Name:
// Module Name: evaluate_network
// Project Name:
// Target Devices:
// Tool Versions:
// Description: Based on Steven's work
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module evaluate_network #(parameter BITS = 16, parameter KERNEL = 7, parameter FEATURES = 21, parameter OVERHEAD_BITS = 12, parameter NB_BASE_BLOCKS = 8, parameter HALF_WIDTH_RAM = 72,
    parameter WIDTH_WEIGHT = 4, parameter WIDTH_FIRST_SIX = 3, parameter WIDTH_OTHERS = 14, parameter BITS_ADDRESS_WEIGHTS = 14, parameter BITS_ADDRESS_BIASES = 9, parameter BITS_ADDRESS_FIRST_SIX = 10,
    parameter BITS_ADDRESS_OTHERS = 12, parameter HALF_CHANNELS_LAYER0 = 4, parameter HALF_CHANNELS_LAYER1 = 16, parameter HALF_CHANNELS_LAYER2 = 32, parameter HALF_CHANNELS_LAYER3 = 16, 
    parameter HALF_CHANNELS_LAYER4 = 8, parameter HALF_CHANNELS_LAYER5 = 1, parameter ROWS_FOR_TILE = 7) (
    input clk,
    input start,
    input [2*BITS-1:0] input_channels,
    input [2:0] stage,
    input [2:0] type,                                               // 000: stage 1, 001: stage 2, 010: left part, 100: middle part, 110: right part. So if third bit is 0 we arrive with 6 clock cycles counter_internal_phase instead of 7. This also applies: layer 5.
    input last_row,
    input [4:0] shift_bias_layer0,
    input [4:0] shift_bias_layer1,
    input [4:0] shift_bias_layer2,
    input [4:0] shift_bias_layer3,
    input [4:0] shift_bias_layer4,
    input [4:0] shift_result_layer0,
    input [4:0] shift_result_layer1,
    input [4:0] shift_result_layer2,
    input [4:0] shift_result_layer3,
    input [4:0] shift_result_layer4,
    output [2*BITS-1:0] output_channels,
    output done
    );

    // Communication with the give_filter_weights block to obtain the filters and biases.
    wire [BITS*KERNEL*NB_BASE_BLOCKS-1:0] filter_weights;
    reg  [BITS*KERNEL*NB_BASE_BLOCKS-1:0] filter_weights_reg = {(BITS*KERNEL*NB_BASE_BLOCKS){1'b0}};
    reg  [2*BITS-1:0] bias_channel = {(2*BITS){1'b0}};
    wire [(2*BITS+OVERHEAD_BITS)*NB_BASE_BLOCKS*KERNEL*(FEATURES-KERNEL+1)-1:0] biases;
    reg  [(2*BITS+OVERHEAD_BITS)*NB_BASE_BLOCKS*KERNEL*(FEATURES-KERNEL+1)-1:0] biases_reg = {(2*BITS+OVERHEAD_BITS)*NB_BASE_BLOCKS*KERNEL*(FEATURES-KERNEL+1){1'b0}};
    reg  [(2*BITS+OVERHEAD_BITS)*4*(FEATURES-KERNEL+1)-1:0] biases_reg_temp_1 = {(2*BITS+OVERHEAD_BITS)*4*(FEATURES-KERNEL+1){1'b0}};
    reg  [(2*BITS+OVERHEAD_BITS)*4*(FEATURES-KERNEL+1)-1:0] biases_reg_temp_2 = {(2*BITS+OVERHEAD_BITS)*4*(FEATURES-KERNEL+1){1'b0}};
    reg  [2*BITS-1:0] output_channels_reg = {(2*BITS){1'b0}};
    reg  [204*(2*BITS+OVERHEAD_BITS)-1:0] results_to_write_in_ram_1 = {(204*(2*BITS+OVERHEAD_BITS)){1'b0}};
    reg  [204*(2*BITS+OVERHEAD_BITS)-1:0] results_to_write_in_ram_2 = {(204*(2*BITS+OVERHEAD_BITS)){1'b0}};
    reg  [2*BITS+OVERHEAD_BITS-1:0] bias_temp1 = {(2*BITS+OVERHEAD_BITS){1'b0}};
    reg  [2*BITS+OVERHEAD_BITS-1:0] bias_temp2 = {(2*BITS+OVERHEAD_BITS){1'b0}};
    assign output_channels = output_channels_reg;
    assign biases = biases_reg;
    assign filter_weights = filter_weights_reg;
    

    // Input and output features for the base blocks
    wire [BITS*NB_BASE_BLOCKS*KERNEL*(FEATURES-KERNEL+1)-1:0] features;
    wire [56*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0] sums1;                 // Not used.
    wire [18*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0] sums3;                 // Not used.
    wire [11*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0] sums5;                 // Not used.
    wire [NB_BASE_BLOCKS*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0] sums7;
    wire [6*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0] sums9;                  // Not used.
    wire [5*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0] sums11;                 // Not used.
    wire [4*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0] sums13;                 // Not used.
    wire [4*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0] results;
   
    
    
    // Counters and help bits for the FSM
    reg  start1 = 1'b1;
    reg  start2 = 1'b0;
    reg  start3 = 1'b0;
    reg  start4 = 1'b0;
    reg  start5 = 1'b0;
    reg  start6 = 1'b0;
    reg  start7 = 1'b0;
    reg  start8 = 1'b0;
    reg  start9 = 1'b0;
    reg  start10 = 1'b0;
    reg  start11 = 1'b0;
    reg  start12 = 1'b0;
    reg  start13 = 1'b0;
    reg  start14 = 1'b0;
    reg  start15 = 1'b0;
    reg  start16 = 1'b0;
    reg  startFSM = 1'b0;
    reg  startUseful = 1'b0;
    reg  start_write_in_ram = 1'b0;
    reg  start_copy_row = 1'b0;
    reg  start_read_new_row = 1'b0;
    reg  start_to_output = 1'b0;
    reg  writing_row = 1'b0;
    reg  continue = 1'b1;
    reg  [15:0] counter_first_phase = {16{1'b0}};           // too many bits, but they still fall away during implementation
    reg  [15:0] counter_internal_phase = {16{1'b0}};
    reg  [15:0] counter_internal_phase_1 = {16{1'b0}};
    reg  [15:0] counter_internal_phase_2 = {16{1'b0}};
    reg  [15:0] counter_internal_phase_3 = {16{1'b0}};
    reg  [15:0] counter_internal_phase_4 = {16{1'b1}};
    reg  [15:0] counter_internal_phase_5 = {16{1'b0}};
    reg  [15:0] counter_internal_phase_6 = {16{1'b0}};
    reg  [15:0] counter_internal_phase_7 = {16{1'b0}};
    reg  [15:0] counter_internal_phase_8 = {16{1'b0}};
    reg  [15:0] counter_internal_phase_9 = {16{1'b0}};
    reg  [15:0] counter_internal_phase_10 = {16{1'b0}};
    reg  [15:0] counterFSM = {16{1'b0}};
    reg  [BITS_ADDRESS_FIRST_SIX-1:0] first_row_data_first_six = {BITS_ADDRESS_FIRST_SIX{1'b0}};
    reg  [BITS_ADDRESS_OTHERS-1:0] first_row_data_others = {BITS_ADDRESS_OTHERS{1'b0}};
    reg  [BITS_ADDRESS_WEIGHTS-1:0] first_row_weights = {BITS_ADDRESS_WEIGHTS{1'b0}};
    reg  [BITS_ADDRESS_BIASES-1:0] first_row_biases = {BITS_ADDRESS_BIASES{1'b0}};
    reg  [BITS_ADDRESS_FIRST_SIX-1:0] first_row_writing_first_six = {BITS_ADDRESS_FIRST_SIX{1'b0}};
    reg  [BITS_ADDRESS_OTHERS-1:0] first_row_writing_others = {BITS_ADDRESS_OTHERS{1'b0}};
    reg  [2:0] row_copy_from = {3{1'b0}};
    reg  [2:0] row_copy_to = {3{1'b0}};
    reg  [6:0] copy_amount_of_channels = 7'b0000000;
    reg  [BITS_ADDRESS_FIRST_SIX-1:0] copy_first_line_first_six = {BITS_ADDRESS_FIRST_SIX{1'b0}};
    reg  [BITS_ADDRESS_OTHERS-1:0] copy_first_line_others = {BITS_ADDRESS_OTHERS{1'b0}};
    reg  [2:0] pointer = {3{1'b0}};
    reg  [2:0] pointer1 = {3{1'b0}};
    reg  [2:0] pointer2 = {3{1'b0}};
    reg  [2:0] pointer3 = {3{1'b0}};
    reg  [2:0] pointer4 = {3{1'b0}};
    reg  [2:0] pointer5 = {3{1'b0}};
    reg  [2:0] layer = {3{1'b0}};
    reg  [5:0] number_two_inputs = 6'b000000;
    reg  [5:0] number_two_outputs = 6'b000000;
    reg  [4:0] shift_bias = {5{1'b0}};
    reg  [4:0] shift_result = {5{1'b0}};
    reg  done_reg = 1'b0;
    assign done = done_reg;
   
    
    // Inputs and outputs of base blocks
    reg  [(2*(FEATURES-KERNEL+1)+(KERNEL-1))*BITS-1:0]   temp_in_1 = {((2*(FEATURES-KERNEL+1)+(KERNEL-1))*BITS){1'b0}};
    reg  [(2*(FEATURES-KERNEL+1)+(KERNEL-1))*BITS-1:0]   temp_in_2 = {((2*(FEATURES-KERNEL+1)+(KERNEL-1))*BITS){1'b0}};
    

    
    
    // Generation of the base_blocks
    base_block_extended #(.BITS(BITS),.OVERHEAD_BITS(OVERHEAD_BITS),.OUTPUTS(FEATURES-KERNEL+1)) base_block_extended(
        .clk(clk),
        .filters(filter_weights),
        .features(features),
        .biases(biases),
        .sums1(sums1),
        .sums3(sums3),
        .sums5(sums5),
        .sums7(sums7),
        .sums9(sums9),
        .sums11(sums11),
        .sums13(sums13)
        );
    genvar ss;
    genvar ww;
    for (ss=0; ss<KERNEL; ss=ss+1)
        begin
            for (ww=0; ww<FEATURES-KERNEL+1; ww=ww+1)
                begin
                    assign features[7*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+(ww+1)*BITS-1:7*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+ww*BITS] = temp_in_1[(FEATURES-KERNEL+1+ss+ww+1)*BITS-1:(FEATURES-KERNEL+1+ss+ww)*BITS];
                    assign features[6*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+(ww+1)*BITS-1:6*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+ww*BITS] = temp_in_2[(FEATURES-KERNEL+1+ss+ww+1)*BITS-1:(FEATURES-KERNEL+1+ss+ww)*BITS];
                    assign features[5*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+(ww+1)*BITS-1:5*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+ww*BITS] = temp_in_1[(ss+ww+1)*BITS-1:(ss+ww)*BITS];
                    assign features[4*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+(ww+1)*BITS-1:4*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+ww*BITS] = temp_in_2[(ss+ww+1)*BITS-1:(ss+ww)*BITS];
                    assign features[3*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+(ww+1)*BITS-1:3*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+ww*BITS] = temp_in_1[(FEATURES-KERNEL+1+ss+ww+1)*BITS-1:(FEATURES-KERNEL+1+ss+ww)*BITS];
                    assign features[2*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+(ww+1)*BITS-1:2*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+ww*BITS] = temp_in_2[(FEATURES-KERNEL+1+ss+ww+1)*BITS-1:(FEATURES-KERNEL+1+ss+ww)*BITS];
                    assign features[1*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+(ww+1)*BITS-1:1*KERNEL*(FEATURES-KERNEL+1)*BITS+ss*(FEATURES-KERNEL+1)*BITS+ww*BITS] = temp_in_1[(ss+ww+1)*BITS-1:(ss+ww)*BITS];
                    assign features[ss*(FEATURES-KERNEL+1)*BITS+(ww+1)*BITS-1:ss*(FEATURES-KERNEL+1)*BITS+ww*BITS] = temp_in_2[(ss+ww+1)*BITS-1:(ss+ww)*BITS];
                end
        end
        
    adder_base_block_extended #(.BITS(BITS),.OVERHEAD_BITS(OVERHEAD_BITS),.NB_BASE_BLOCKS(NB_BASE_BLOCKS), 
    .FEATURES(FEATURES),.KERNEL(KERNEL)) adder_base_block_extended(
            .clk(clk),
            .sums7(sums7),
            .results(results)
            );
    
    
    wire en;
    wire write_weightsOddInputChannelOddOutputChannel;
    wire write_weightsOddInputChannelEvenOutputChannel;
    wire write_weightsEvenInputChannelOddOutputChannel;
    wire write_weightsEvenInputChannelEvenOutputChannel;
    wire write_biasesMemory;
    wire write_firstWordsOddChannels;
    wire write_firstWordsEvenChannels;
    wire write_otherWordsOddChannels;
    wire write_otherWordsEvenChannels;
    wire [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsOddInputChannelOddOutputChannel_input;
    wire [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsOddInputChannelEvenOutputChannel_input;
    wire [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsEvenInputChannelOddOutputChannel_input;
    wire [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsEvenInputChannelEvenOutputChannel_input;
    wire [HALF_WIDTH_RAM-1:0] biasesMemory_input;
    wire [HALF_WIDTH_RAM*WIDTH_FIRST_SIX-1:0] firstWordsOddChannels_input;
    wire [HALF_WIDTH_RAM*WIDTH_FIRST_SIX-1:0] firstWordsEvenChannels_input;
    wire [HALF_WIDTH_RAM*WIDTH_OTHERS-1:0] otherWordsOddChannels_input;
    wire [HALF_WIDTH_RAM*WIDTH_OTHERS-1:0] otherWordsEvenChannels_input;
    wire [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsOddInputChannelOddOutputChannel_output;
    wire [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsOddInputChannelEvenOutputChannel_output;
    wire [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsEvenInputChannelOddOutputChannel_output;
    wire [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsEvenInputChannelEvenOutputChannel_output;
    wire [HALF_WIDTH_RAM-1:0] biasesMemory_output;
    wire [HALF_WIDTH_RAM*WIDTH_FIRST_SIX-1:0] firstWordsOddChannels_output;
    wire [HALF_WIDTH_RAM*WIDTH_FIRST_SIX-1:0] firstWordsEvenChannels_output;
    wire [HALF_WIDTH_RAM*WIDTH_OTHERS-1:0] otherWordsOddChannels_output; 
    wire [HALF_WIDTH_RAM*WIDTH_OTHERS-1:0] otherWordsEvenChannels_output;
    wire [BITS_ADDRESS_WEIGHTS-1:0] read_address_weightsOddInputChannelOddOutputChannel;
    wire [BITS_ADDRESS_WEIGHTS-1:0] read_address_weightsOddInputChannelEvenOutputChannel;
    wire [BITS_ADDRESS_WEIGHTS-1:0] read_address_weightsEvenInputChannelOddOutputChannel;
    wire [BITS_ADDRESS_WEIGHTS-1:0] read_address_weightsEvenInputChannelEvenOutputChannel;
    wire [BITS_ADDRESS_BIASES-1:0] read_address_biasesMemory;
    wire [BITS_ADDRESS_FIRST_SIX-1:0] read_address_firstWordsOddChannels;
    wire [BITS_ADDRESS_FIRST_SIX-1:0] read_address_firstWordsEvenChannels;
    wire [BITS_ADDRESS_OTHERS-1:0] read_address_otherWordsOddChannels;
    wire [BITS_ADDRESS_OTHERS-1:0] read_address_otherWordsEvenChannels;
    wire [BITS_ADDRESS_WEIGHTS-1:0] write_address_weightsOddInputChannelOddOutputChannel;
    wire [BITS_ADDRESS_WEIGHTS-1:0] write_address_weightsOddInputChannelEvenOutputChannel;
    wire [BITS_ADDRESS_WEIGHTS-1:0] write_address_weightsEvenInputChannelOddOutputChannel;
    wire [BITS_ADDRESS_WEIGHTS-1:0] write_address_weightsEvenInputChannelEvenOutputChannel;
    wire [BITS_ADDRESS_BIASES-1:0] write_address_biasesMemory;
    wire [BITS_ADDRESS_FIRST_SIX-1:0] write_address_firstWordsOddChannels;
    wire [BITS_ADDRESS_FIRST_SIX-1:0] write_address_firstWordsEvenChannels;
    wire [BITS_ADDRESS_OTHERS-1:0] write_address_otherWordsOddChannels;
    wire [BITS_ADDRESS_OTHERS-1:0] write_address_otherWordsEvenChannels;
    reg  en_reg = 1'b1;
    reg  write_weightsOddInputChannelOddOutputChannel_reg = 1'b0;
    reg  write_weightsOddInputChannelEvenOutputChannel_reg = 1'b0;
    reg  write_weightsEvenInputChannelOddOutputChannel_reg = 1'b0;
    reg  write_weightsEvenInputChannelEvenOutputChannel_reg = 1'b0;
    reg  write_biasesMemory_reg = 1'b0;
    reg  write_firstWordsOddChannels_reg = 1'b0;
    reg  write_firstWordsEvenChannels_reg = 1'b0;
    reg  write_otherWordsOddChannels_reg = 1'b0; 
    reg  write_otherWordsEvenChannels_reg = 1'b0;
    reg [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsOddInputChannelOddOutputChannel_input_reg = {(HALF_WIDTH_RAM*WIDTH_WEIGHT){1'b0}};
    reg [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsOddInputChannelEvenOutputChannel_input_reg = {(HALF_WIDTH_RAM*WIDTH_WEIGHT){1'b0}};
    reg [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsEvenInputChannelOddOutputChannel_input_reg = {(HALF_WIDTH_RAM*WIDTH_WEIGHT){1'b0}};
    reg [HALF_WIDTH_RAM*WIDTH_WEIGHT-1:0] weightsEvenInputChannelEvenOutputChannel_input_reg = {(HALF_WIDTH_RAM*WIDTH_WEIGHT){1'b0}};
    reg [HALF_WIDTH_RAM-1:0] biasesMemory_input_reg = {(HALF_WIDTH_RAM){1'b0}};
    reg [HALF_WIDTH_RAM*WIDTH_FIRST_SIX-1:0] firstWordsOddChannels_input_reg = {(HALF_WIDTH_RAM*WIDTH_FIRST_SIX){1'b0}};
    reg [HALF_WIDTH_RAM*WIDTH_FIRST_SIX-1:0] firstWordsEvenChannels_input_reg = {(HALF_WIDTH_RAM*WIDTH_FIRST_SIX){1'b0}};
    reg [HALF_WIDTH_RAM*WIDTH_OTHERS-1:0] otherWordsOddChannels_input_reg = {(HALF_WIDTH_RAM*WIDTH_OTHERS){1'b0}}; 
    reg [HALF_WIDTH_RAM*WIDTH_OTHERS-1:0] otherWordsEvenChannels_input_reg = {(HALF_WIDTH_RAM*WIDTH_OTHERS){1'b0}};
    reg [BITS_ADDRESS_WEIGHTS-1:0] read_address_weightsOddInputChannelOddOutputChannel_reg = {BITS_ADDRESS_WEIGHTS{1'b0}};
    reg [BITS_ADDRESS_WEIGHTS-1:0] read_address_weightsOddInputChannelEvenOutputChannel_reg = {BITS_ADDRESS_WEIGHTS{1'b0}};
    reg [BITS_ADDRESS_WEIGHTS-1:0] read_address_weightsEvenInputChannelOddOutputChannel_reg = {BITS_ADDRESS_WEIGHTS{1'b0}};
    reg [BITS_ADDRESS_WEIGHTS-1:0] read_address_weightsEvenInputChannelEvenOutputChannel_reg = {BITS_ADDRESS_WEIGHTS{1'b0}};
    reg [BITS_ADDRESS_BIASES-1:0] read_address_biasesMemory_reg = {BITS_ADDRESS_BIASES{1'b0}};
    reg [BITS_ADDRESS_FIRST_SIX-1:0] read_address_firstWordsOddChannels_reg = {BITS_ADDRESS_FIRST_SIX{1'b0}};
    reg [BITS_ADDRESS_FIRST_SIX-1:0] read_address_firstWordsEvenChannels_reg = {BITS_ADDRESS_FIRST_SIX{1'b0}};
    reg [BITS_ADDRESS_OTHERS-1:0] read_address_otherWordsOddChannels_reg = {BITS_ADDRESS_OTHERS{1'b0}};
    reg [BITS_ADDRESS_OTHERS-1:0] read_address_otherWordsEvenChannels_reg = {BITS_ADDRESS_OTHERS{1'b0}};
    reg [BITS_ADDRESS_WEIGHTS-1:0] write_address_weightsOddInputChannelOddOutputChannel_reg = {BITS_ADDRESS_WEIGHTS{1'b0}};
    reg [BITS_ADDRESS_WEIGHTS-1:0] write_address_weightsOddInputChannelEvenOutputChannel_reg = {BITS_ADDRESS_WEIGHTS{1'b0}};
    reg [BITS_ADDRESS_WEIGHTS-1:0] write_address_weightsEvenInputChannelOddOutputChannel_reg = {BITS_ADDRESS_WEIGHTS{1'b0}};
    reg [BITS_ADDRESS_WEIGHTS-1:0] write_address_weightsEvenInputChannelEvenOutputChannel_reg = {BITS_ADDRESS_WEIGHTS{1'b0}};
    reg [BITS_ADDRESS_BIASES-1:0] write_address_biasesMemory_reg = {BITS_ADDRESS_BIASES{1'b0}};
    reg [BITS_ADDRESS_FIRST_SIX-1:0] write_address_firstWordsOddChannels_reg = {BITS_ADDRESS_FIRST_SIX{1'b0}};
    reg [BITS_ADDRESS_FIRST_SIX-1:0] write_address_firstWordsEvenChannels_reg = {BITS_ADDRESS_FIRST_SIX{1'b0}};
    reg [BITS_ADDRESS_OTHERS-1:0] write_address_otherWordsOddChannels_reg = {BITS_ADDRESS_OTHERS{1'b0}};
    reg [BITS_ADDRESS_OTHERS-1:0] write_address_otherWordsEvenChannels_reg = {BITS_ADDRESS_OTHERS{1'b0}};
    assign en = en_reg;
    assign write_weightsOddInputChannelOddOutputChannel = write_weightsOddInputChannelOddOutputChannel_reg;
    assign write_weightsOddInputChannelEvenOutputChannel = write_weightsOddInputChannelEvenOutputChannel_reg;
    assign write_weightsEvenInputChannelOddOutputChannel = write_weightsEvenInputChannelOddOutputChannel_reg;
    assign write_weightsEvenInputChannelEvenOutputChannel = write_weightsEvenInputChannelEvenOutputChannel_reg;
    assign write_biasesMemory = write_biasesMemory_reg;
    assign write_firstWordsOddChannels = write_firstWordsOddChannels_reg;
    assign write_firstWordsEvenChannels = write_firstWordsEvenChannels_reg;
    assign write_otherWordsOddChannels = write_otherWordsOddChannels_reg;
    assign write_otherWordsEvenChannels = write_otherWordsEvenChannels_reg;
    assign weightsOddInputChannelOddOutputChannel_input = weightsOddInputChannelOddOutputChannel_input_reg;
    assign weightsOddInputChannelEvenOutputChannel_input = weightsOddInputChannelEvenOutputChannel_input_reg;
    assign weightsEvenInputChannelOddOutputChannel_input = weightsEvenInputChannelOddOutputChannel_input_reg;
    assign weightsEvenInputChannelEvenOutputChannel_input = weightsEvenInputChannelEvenOutputChannel_input_reg;
    assign biasesMemory_input = biasesMemory_input_reg;
    assign firstWordsOddChannels_input = firstWordsOddChannels_input_reg;
    assign firstWordsEvenChannels_input = firstWordsEvenChannels_input_reg;
    assign otherWordsOddChannels_input = otherWordsOddChannels_input_reg;
    assign otherWordsEvenChannels_input = otherWordsEvenChannels_input_reg;
    assign read_address_weightsOddInputChannelOddOutputChannel = read_address_weightsOddInputChannelOddOutputChannel_reg;
    assign read_address_weightsOddInputChannelEvenOutputChannel = read_address_weightsOddInputChannelEvenOutputChannel_reg;
    assign read_address_weightsEvenInputChannelOddOutputChannel = read_address_weightsEvenInputChannelOddOutputChannel_reg;
    assign read_address_weightsEvenInputChannelEvenOutputChannel = read_address_weightsEvenInputChannelEvenOutputChannel_reg;
    assign read_address_biasesMemory = read_address_biasesMemory_reg;
    assign read_address_firstWordsOddChannels = read_address_firstWordsOddChannels_reg;
    assign read_address_firstWordsEvenChannels = read_address_firstWordsEvenChannels_reg;
    assign read_address_otherWordsOddChannels = read_address_otherWordsOddChannels_reg;
    assign read_address_otherWordsEvenChannels = read_address_otherWordsEvenChannels_reg;
    assign write_address_weightsOddInputChannelOddOutputChannel = write_address_weightsOddInputChannelOddOutputChannel_reg;
    assign write_address_weightsOddInputChannelEvenOutputChannel = write_address_weightsOddInputChannelEvenOutputChannel_reg;
    assign write_address_weightsEvenInputChannelOddOutputChannel = write_address_weightsEvenInputChannelOddOutputChannel_reg;
    assign write_address_weightsEvenInputChannelEvenOutputChannel = write_address_weightsEvenInputChannelEvenOutputChannel_reg;
    assign write_address_biasesMemory = write_address_biasesMemory_reg;
    assign write_address_firstWordsOddChannels = write_address_firstWordsOddChannels_reg;
    assign write_address_firstWordsEvenChannels = write_address_firstWordsEvenChannels_reg;
    assign write_address_otherWordsOddChannels = write_address_otherWordsOddChannels_reg;
    assign write_address_otherWordsEvenChannels = write_address_otherWordsEvenChannels_reg;
    //
    blk_mem_gen_2 weightsOddInputChannelOddOutputChannel (
          .clka(clk),    
          .ena(en),      
          .wea(write_weightsOddInputChannelOddOutputChannel),      
          .addra(write_address_weightsOddInputChannelOddOutputChannel),  
          .dina(weightsOddInputChannelOddOutputChannel_input),    
          .clkb(clk),   
          .enb(en),      
          .addrb(read_address_weightsOddInputChannelOddOutputChannel),  
          .doutb(weightsOddInputChannelOddOutputChannel_output)  
        );
    blk_mem_gen_2 weightsOddInputChannelEvenOutputChannel (
          .clka(clk),    
          .ena(en),      
          .wea(write_weightsOddInputChannelEvenOutputChannel),     
          .addra(write_address_weightsOddInputChannelEvenOutputChannel),  
          .dina(weightsOddInputChannelEvenOutputChannel_input),    
          .clkb(clk),    
          .enb(en),      
          .addrb(read_address_weightsOddInputChannelEvenOutputChannel),  
          .doutb(weightsOddInputChannelEvenOutputChannel_output)  
        );
    blk_mem_gen_2 weightsEvenInputChannelOddOutputChannel (
          .clka(clk),    
          .ena(en),      
          .wea(write_weightsEvenInputChannelOddOutputChannel),      
          .addra(write_address_weightsEvenInputChannelOddOutputChannel),  
          .dina(weightsEvenInputChannelOddOutputChannel_input),    
          .clkb(clk),    
          .enb(en),     
          .addrb(read_address_weightsEvenInputChannelOddOutputChannel),  
          .doutb(weightsEvenInputChannelOddOutputChannel_output) 
        );
    blk_mem_gen_2 weightsEvenInputChannelEvenOutputChannel (
          .clka(clk),    
          .ena(en),     
          .wea(write_weightsEvenInputChannelEvenOutputChannel),      
          .addra(write_address_weightsEvenInputChannelEvenOutputChannel),  
          .dina(weightsEvenInputChannelEvenOutputChannel_input),   
          .clkb(clk),    
          .enb(en),      
          .addrb(read_address_weightsEvenInputChannelEvenOutputChannel),  
          .doutb(weightsEvenInputChannelEvenOutputChannel_output)
        );
    blk_mem_gen_1 biasesMemory (
          .clka(clk),   
          .ena(en),      
          .wea(write_biasesMemory),      
          .addra(write_address_biasesMemory),  
          .dina(biasesMemory_input),   
          .clkb(clk),    
          .enb(en),      
          .addrb(read_address_biasesMemory),  
          .doutb(biasesMemory_output)  
        );
    blk_mem_gen_3 firstWordsOddChannels (
          .clka(clk),    
          .ena(en),      
          .wea(write_firstWordsOddChannels),      
          .addra(write_address_firstWordsOddChannels),  
          .dina(firstWordsOddChannels_input),    
          .clkb(clk),  
          .enb(en),    
          .addrb(read_address_firstWordsOddChannels),  
          .doutb(firstWordsOddChannels_output)  
        );
    blk_mem_gen_3 firstWordsEvenChannels (
          .clka(clk),   
          .ena(en),      
          .wea(write_firstWordsEvenChannels),     
          .addra(write_address_firstWordsEvenChannels),  
          .dina(firstWordsEvenChannels_input),    
          .clkb(clk),    
          .enb(en),      
          .addrb(read_address_firstWordsEvenChannels),  
          .doutb(firstWordsEvenChannels_output)  
        );
    blk_mem_gen_4 otherWordsOddChannels (
          .clka(clk),    
          .ena(en),      
          .wea(write_otherWordsOddChannels),      
          .addra(write_address_otherWordsOddChannels),  
          .dina(otherWordsOddChannels_input),    
          .clkb(clk),  
          .enb(en),    
          .addrb(read_address_otherWordsOddChannels),  
          .doutb(otherWordsOddChannels_output)  
        );
    blk_mem_gen_4 otherWordsEvenChannels (
          .clka(clk),   
          .ena(en),      
          .wea(write_otherWordsEvenChannels),     
          .addra(write_address_otherWordsEvenChannels),  
          .dina(otherWordsEvenChannels_input),    
          .clkb(clk),    
          .enb(en),      
          .addrb(read_address_otherWordsEvenChannels),  
          .doutb(otherWordsEvenChannels_output)  
        );
    always @(posedge clk)
    begin
    if (start == 1)
        begin
            if (start1 == 1) 
                begin
                    case(counter_first_phase)
                    1   :   weightsOddInputChannelOddOutputChannel_input_reg[7*BITS-1:5*BITS] <= input_channels;
                    2   :   weightsOddInputChannelOddOutputChannel_input_reg[5*BITS-1:3*BITS] <= input_channels;
                    3   :   weightsOddInputChannelOddOutputChannel_input_reg[3*BITS-1:BITS] <= input_channels;
                    0   :   weightsOddInputChannelOddOutputChannel_input_reg[BITS-1:0] <= input_channels[2*BITS-1:BITS];
                    endcase
                    if (counter_first_phase == 3)
                        begin
                            counter_first_phase <= 0;
                            if (counter_internal_phase_1 == KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + 
                                HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4 + HALF_CHANNELS_LAYER4*HALF_CHANNELS_LAYER5) - 1)
                                begin
                                start1 <= 0;
                                start2 <= 1;
                                counter_internal_phase_1 <= 0;
                                end
                            else
                                counter_internal_phase_1 <= counter_internal_phase_1 + 1;
                        end
                    else if (counter_first_phase == 0)
                        begin
                            counter_first_phase <= counter_first_phase + 1;
                            write_weightsOddInputChannelOddOutputChannel_reg <= 1;
                            if (counter_internal_phase_1 != 0)
                                write_address_weightsOddInputChannelOddOutputChannel_reg <= counter_internal_phase_1 - 1;
                        end
                    else
                        begin
                            counter_first_phase <= counter_first_phase + 1;
                            write_weightsOddInputChannelOddOutputChannel_reg <= 0;
                        end
                end
        end
    else
        begin
            start1 <= 1;
        end
    if (start2 == 1)
        begin
            case(counter_first_phase)
            1   :   weightsOddInputChannelEvenOutputChannel_input_reg[7*BITS-1:5*BITS] <= input_channels;
            2   :   weightsOddInputChannelEvenOutputChannel_input_reg[5*BITS-1:3*BITS] <= input_channels;
            3   :   weightsOddInputChannelEvenOutputChannel_input_reg[3*BITS-1:BITS] <= input_channels;
            0   :   weightsOddInputChannelEvenOutputChannel_input_reg[BITS-1:0] <= input_channels[2*BITS-1:BITS];
            endcase
            if (counter_first_phase == 3)
                begin
                    counter_first_phase <= 0;
                    if (counter_internal_phase_1 == KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + 
                        HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4 + HALF_CHANNELS_LAYER4*HALF_CHANNELS_LAYER5) - 1)
                        begin
                        start2 <= 0;
                        start3 <= 1;
                        counter_internal_phase_1 <= 0;
                        end
                    else
                        counter_internal_phase_1 <= counter_internal_phase_1 + 1;
                end
            else if (counter_first_phase == 0)
                begin
                counter_first_phase <= counter_first_phase + 1;
                    if (counter_internal_phase_1 == 0)
                        begin
                        write_weightsOddInputChannelOddOutputChannel_reg <= 1;
                        write_address_weightsOddInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + 
                        HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4 + HALF_CHANNELS_LAYER4*HALF_CHANNELS_LAYER5) - 1;
                        end
                    else
                        begin
                        write_weightsOddInputChannelEvenOutputChannel_reg <= 1;
                        write_address_weightsOddInputChannelEvenOutputChannel_reg <= counter_internal_phase_1 - 1;
                        end
                    end
            else 
                begin
                    write_weightsOddInputChannelOddOutputChannel_reg <= 0;
                    write_weightsOddInputChannelEvenOutputChannel_reg <= 0;
                    counter_first_phase <= counter_first_phase + 1;
                end
        end
    if (start3 == 1)
            begin
                case(counter_first_phase)
                1   :   weightsEvenInputChannelOddOutputChannel_input_reg[7*BITS-1:5*BITS] <= input_channels;
                2   :   weightsEvenInputChannelOddOutputChannel_input_reg[5*BITS-1:3*BITS] <= input_channels;
                3   :   weightsEvenInputChannelOddOutputChannel_input_reg[3*BITS-1:BITS] <= input_channels;
                0   :   weightsEvenInputChannelOddOutputChannel_input_reg[BITS-1:0] <= input_channels[2*BITS-1:BITS];
                endcase
                if (counter_first_phase == 3)
                    begin
                        counter_first_phase <= 0;
                        if (counter_internal_phase_1 == KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + 
                            HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4 + HALF_CHANNELS_LAYER4*HALF_CHANNELS_LAYER5) - 1)
                            begin
                            start3 <= 0;
                            start4 <= 1;
                            counter_internal_phase_1 <= 0;
                            end
                        else
                            counter_internal_phase_1 <= counter_internal_phase_1 + 1;
                    end
                else if (counter_first_phase == 0)
                    begin
                    counter_first_phase <= counter_first_phase + 1;
                        if (counter_internal_phase_1 == 0)
                            begin
                            write_weightsOddInputChannelEvenOutputChannel_reg <= 1;
                            write_address_weightsOddInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + 
                            HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4 + HALF_CHANNELS_LAYER4*HALF_CHANNELS_LAYER5)- 1;
                            end
                        else
                            begin
                            write_weightsEvenInputChannelOddOutputChannel_reg <= 1;
                            write_address_weightsEvenInputChannelOddOutputChannel_reg <= counter_internal_phase_1 - 1;
                            end
                        end
                else 
                    begin
                        write_weightsOddInputChannelEvenOutputChannel_reg <= 0;
                        write_weightsEvenInputChannelOddOutputChannel_reg <= 0;
                        counter_first_phase <= counter_first_phase + 1;
                    end
            end
     if (start4 == 1)
            begin
                case(counter_first_phase)
                1   :   weightsEvenInputChannelEvenOutputChannel_input_reg[7*BITS-1:5*BITS] <= input_channels;
                2   :   weightsEvenInputChannelEvenOutputChannel_input_reg[5*BITS-1:3*BITS] <= input_channels;
                3   :   weightsEvenInputChannelEvenOutputChannel_input_reg[3*BITS-1:BITS] <= input_channels;
                0   :   weightsEvenInputChannelEvenOutputChannel_input_reg[BITS-1:0] <= input_channels[2*BITS-1:BITS];
                endcase
                if (counter_first_phase == 3)
                    begin
                        counter_first_phase <= 0;
                        if (counter_internal_phase_1 == KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + 
                            HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4 + HALF_CHANNELS_LAYER4*HALF_CHANNELS_LAYER5) - 1)
                            begin
                            start4 <= 0;
                            start5 <= 1;
                            counter_internal_phase_1 <= 0;
                            end
                        else
                            counter_internal_phase_1 <= counter_internal_phase_1 + 1;
                    end
                else if (counter_first_phase == 0)
                    begin
                    counter_first_phase <= counter_first_phase + 1;
                        if (counter_internal_phase_1 == 0)
                            begin
                            write_weightsEvenInputChannelOddOutputChannel_reg <= 1;
                            write_address_weightsEvenInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + 
                            HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4 + HALF_CHANNELS_LAYER4*HALF_CHANNELS_LAYER5) - 1;
                            end
                        else
                            begin
                            write_weightsEvenInputChannelEvenOutputChannel_reg <= 1;
                            write_address_weightsEvenInputChannelEvenOutputChannel_reg <= counter_internal_phase_1 - 1;
                            end
                        end
                else 
                    begin
                        write_weightsEvenInputChannelEvenOutputChannel_reg <= 0;
                        write_weightsEvenInputChannelOddOutputChannel_reg <= 0;
                        counter_first_phase <= counter_first_phase + 1;
                    end
            end
    if (start5 == 1)
        begin
            if (counter_first_phase == 0)
                begin
                counter_first_phase <= counter_first_phase + 1;
                weightsEvenInputChannelEvenOutputChannel_input_reg[BITS-1:0] <= input_channels[2*BITS-1:BITS];
                write_weightsEvenInputChannelEvenOutputChannel_reg <= 1;
                write_address_weightsEvenInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + 
                HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4 + HALF_CHANNELS_LAYER4*HALF_CHANNELS_LAYER5) - 1;
                end
            else 
                begin
                biasesMemory_input_reg[2*BITS-1:0] <= input_channels;
                write_weightsEvenInputChannelEvenOutputChannel_reg <= 0;
                write_biasesMemory_reg <= 1;
                write_address_biasesMemory_reg <= counter_first_phase - 1;
                if (counter_first_phase == HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER4 + HALF_CHANNELS_LAYER5)
                    begin
                    start5 <= 0;
                    start6 <= 1;
                    counter_first_phase <= 0;
                    counter_internal_phase_1 <= 0;
                    end
                else
                    counter_first_phase <= counter_first_phase + 1;
                end
        end   
    if (start6 == 1)   
        begin
        write_biasesMemory_reg <= 0;
        case(counter_first_phase)
        0   :   firstWordsOddChannels_input_reg[6*BITS-1:4*BITS] <= input_channels;
        1   :   firstWordsOddChannels_input_reg[4*BITS-1:2*BITS] <= input_channels;
        2   :   firstWordsOddChannels_input_reg[2*BITS-1:0] <= input_channels;
        endcase
        if (counter_first_phase == 2)
            begin
                counter_first_phase <= 0;
                write_firstWordsOddChannels_reg <= 1;
                write_address_firstWordsOddChannels_reg <= KERNEL*counter_internal_phase_1[10:2] + 3 + counter_internal_phase_1[1:0];
                if (counter_internal_phase_1 == 4*HALF_CHANNELS_LAYER0 - 1)
                    begin
                    start6 <= 0;
                    start7 <= 1;
                    counter_internal_phase_1 <= 0;
                    end
                else
                    counter_internal_phase_1 <= counter_internal_phase_1 + 1;
            end
        else 
            begin
                write_firstWordsOddChannels_reg <= 0;
                counter_first_phase <= counter_first_phase + 1;
            end
        end
    if (start7 == 1)   
        begin
        write_firstWordsOddChannels_reg <= 0;
        case(counter_first_phase)
        0   :   firstWordsEvenChannels_input_reg[6*BITS-1:4*BITS] <= input_channels;
        1   :   firstWordsEvenChannels_input_reg[4*BITS-1:2*BITS] <= input_channels;
        2   :   firstWordsEvenChannels_input_reg[2*BITS-1:0] <= input_channels;
        endcase
        if (counter_first_phase == 2)
            begin
                counter_first_phase <= 0;
                write_firstWordsEvenChannels_reg <= 1;
                write_address_firstWordsEvenChannels_reg <= KERNEL*counter_internal_phase_1[10:2] + 3 + counter_internal_phase_1[1:0];
                if (counter_internal_phase_1 == 4*HALF_CHANNELS_LAYER0 - 1)
                    begin
                    start7 <= 0;
                    start8 <= 1;
                    counter_internal_phase_1 <= 0;
                    counter_internal_phase <= 0;
                    end
                else
                    counter_internal_phase_1 <= counter_internal_phase_1 + 1;
            end
        else 
            begin
                write_firstWordsEvenChannels_reg <= 0;
                counter_first_phase <= counter_first_phase + 1;
            end
        end
    if (start8 == 1)   
        begin
        write_firstWordsEvenChannels_reg <= 0;
        case(counter_first_phase)
        0   :   otherWordsOddChannels_input_reg[30*BITS-1:28*BITS] <= input_channels;
        1   :   otherWordsOddChannels_input_reg[28*BITS-1:26*BITS] <= input_channels;
        2   :   otherWordsOddChannels_input_reg[26*BITS-1:24*BITS] <= input_channels;
        3   :   otherWordsOddChannels_input_reg[24*BITS-1:22*BITS] <= input_channels;
        4   :   otherWordsOddChannels_input_reg[22*BITS-1:20*BITS] <= input_channels;
        5   :   otherWordsOddChannels_input_reg[20*BITS-1:18*BITS] <= input_channels;
        6   :   otherWordsOddChannels_input_reg[18*BITS-1:16*BITS] <= input_channels;
        7   :   otherWordsOddChannels_input_reg[16*BITS-1:14*BITS] <= input_channels;
        8   :   otherWordsOddChannels_input_reg[14*BITS-1:12*BITS] <= input_channels;
        9   :   otherWordsOddChannels_input_reg[12*BITS-1:10*BITS] <= input_channels;
        10   :   otherWordsOddChannels_input_reg[10*BITS-1:8*BITS] <= input_channels;
        11   :   otherWordsOddChannels_input_reg[8*BITS-1:6*BITS] <= input_channels;
        12   :   otherWordsOddChannels_input_reg[6*BITS-1:4*BITS] <= input_channels;
        13   :   otherWordsOddChannels_input_reg[4*BITS-1:2*BITS] <= input_channels;
        14   :   otherWordsOddChannels_input_reg[2*BITS-1:0] <= input_channels;
        endcase
        if (counter_first_phase == 14)
            begin
                counter_first_phase <= 0;
                write_otherWordsOddChannels_reg <= 1;
                write_address_otherWordsOddChannels_reg <= KERNEL*ROWS_FOR_TILE*counter_internal_phase_1[10:2] + ROWS_FOR_TILE*(3+counter_internal_phase_1[1:0]) + counter_internal_phase;
                if (counter_internal_phase_1 == 4*HALF_CHANNELS_LAYER0 - 1)
                    if (counter_internal_phase == ROWS_FOR_TILE - 1)
                        begin
                        start8 <= 0;
                        start9 <= 1;
                        counter_internal_phase_1 <= 0;
                        counter_internal_phase <= 0;
                        end
                    else
                        counter_internal_phase <= counter_internal_phase + 1;
                else
                    begin
                    if (counter_internal_phase == ROWS_FOR_TILE - 1)
                        begin
                            counter_internal_phase_1 <= counter_internal_phase_1 + 1;
                            counter_internal_phase <= 0;
                        end
                    else
                        counter_internal_phase <= counter_internal_phase + 1;
                    end
            end
        else 
            begin
                write_otherWordsOddChannels_reg <= 0;
                counter_first_phase <= counter_first_phase + 1;
            end
        end
    if (start9 == 1)   
        begin
        write_otherWordsOddChannels_reg <= 0;
        case(counter_first_phase)
        0   :   otherWordsEvenChannels_input_reg[30*BITS-1:28*BITS] <= input_channels;
        1   :   otherWordsEvenChannels_input_reg[28*BITS-1:26*BITS] <= input_channels;
        2   :   otherWordsEvenChannels_input_reg[26*BITS-1:24*BITS] <= input_channels;
        3   :   otherWordsEvenChannels_input_reg[24*BITS-1:22*BITS] <= input_channels;
        4   :   otherWordsEvenChannels_input_reg[22*BITS-1:20*BITS] <= input_channels;
        5   :   otherWordsEvenChannels_input_reg[20*BITS-1:18*BITS] <= input_channels;
        6   :   otherWordsEvenChannels_input_reg[18*BITS-1:16*BITS] <= input_channels;
        7   :   otherWordsEvenChannels_input_reg[16*BITS-1:14*BITS] <= input_channels;
        8   :   otherWordsEvenChannels_input_reg[14*BITS-1:12*BITS] <= input_channels;
        9   :   otherWordsEvenChannels_input_reg[12*BITS-1:10*BITS] <= input_channels;
        10   :   otherWordsEvenChannels_input_reg[10*BITS-1:8*BITS] <= input_channels;
        11   :   otherWordsEvenChannels_input_reg[8*BITS-1:6*BITS] <= input_channels;
        12   :   otherWordsEvenChannels_input_reg[6*BITS-1:4*BITS] <= input_channels;
        13   :   otherWordsEvenChannels_input_reg[4*BITS-1:2*BITS] <= input_channels;
        14   :   otherWordsEvenChannels_input_reg[2*BITS-1:0] <= input_channels;
        endcase
        if (counter_first_phase == 14)
            begin
                counter_first_phase <= 0;
                write_otherWordsEvenChannels_reg <= 1;
                write_address_otherWordsEvenChannels_reg <= KERNEL*ROWS_FOR_TILE*counter_internal_phase_1[10:2] + ROWS_FOR_TILE*(3+counter_internal_phase_1[1:0]) + counter_internal_phase;
                if (counter_internal_phase_1 == 4*HALF_CHANNELS_LAYER0 - 1)
                    if (counter_internal_phase == ROWS_FOR_TILE - 1)
                        begin
                        start9 <= 0;
                        start10 <= 1;
                        counter_internal_phase_1 <= 0;
                        counter_internal_phase <= 0;
                        end
                    else
                        counter_internal_phase <= counter_internal_phase + 1;
                else
                    begin
                    if (counter_internal_phase == ROWS_FOR_TILE - 1)
                        begin
                            counter_internal_phase_1 <= counter_internal_phase_1 + 1;
                            counter_internal_phase <= 0;
                        end
                    else
                        counter_internal_phase <= counter_internal_phase + 1;
                    end
            end
        else 
            begin
                write_otherWordsEvenChannels_reg <= 0;
                counter_first_phase <= counter_first_phase + 1;
            end
        end
    if (start_copy_row == 1)
        begin
        otherWordsOddChannels_input_reg[2*(FEATURES-KERNEL+1)*BITS-1:0] <= otherWordsOddChannels_output[2*(FEATURES-KERNEL+1)*BITS-1:0];
        otherWordsEvenChannels_input_reg[2*(FEATURES-KERNEL+1)*BITS-1:0] <= otherWordsEvenChannels_output[2*(FEATURES-KERNEL+1)*BITS-1:0];
        firstWordsOddChannels_input_reg[(KERNEL-1)*BITS-1:0] <= firstWordsOddChannels_output[(KERNEL-1)*BITS-1:0];
        firstWordsEvenChannels_input_reg[(KERNEL-1)*BITS-1:0] <= firstWordsEvenChannels_output[(KERNEL-1)*BITS-1:0];
        if (counter_internal_phase_7 != copy_amount_of_channels)
            begin
                read_address_otherWordsOddChannels_reg <= copy_first_line_others + ROWS_FOR_TILE*row_copy_from + KERNEL*ROWS_FOR_TILE*counter_internal_phase_7 + counter_internal_phase_8;
                read_address_otherWordsEvenChannels_reg <= copy_first_line_others + ROWS_FOR_TILE*row_copy_from + KERNEL*ROWS_FOR_TILE*counter_internal_phase_7 + counter_internal_phase_8;
                read_address_firstWordsOddChannels_reg <= copy_first_line_first_six + row_copy_from + KERNEL*counter_internal_phase_7;
                read_address_firstWordsEvenChannels_reg <= copy_first_line_first_six + row_copy_from + KERNEL*counter_internal_phase_7;
            end
        if (counter_internal_phase_8 == ROWS_FOR_TILE-1)
            begin
            counter_internal_phase_8 <= 0;
            counter_internal_phase_7 <= counter_internal_phase_7 + 1;
            end
        else
            begin
            counter_internal_phase_8 <= counter_internal_phase_8 + 1;
            if (counter_internal_phase_8 == 3)  
                begin
                if (counter_internal_phase_7 == copy_amount_of_channels)
                    begin
                    start_copy_row <= 0;
                    counter_internal_phase_7 <= 0;
                    counter_internal_phase_8 <= 0;
                    write_otherWordsOddChannels_reg <= 0;
                    write_otherWordsEvenChannels_reg <= 0;
                    end
                else
                    begin
                    write_otherWordsOddChannels_reg <= 1;
                    write_otherWordsEvenChannels_reg <= 1;
                    write_firstWordsOddChannels_reg <= 1;
                    write_firstWordsEvenChannels_reg <= 1;
                    end
                end
            if (counter_internal_phase_8 == 4)
                begin
                write_firstWordsOddChannels_reg <= 0;
                write_firstWordsEvenChannels_reg <= 0;
                end
            end
        if (counter_internal_phase_8 >= 3)
            begin
            write_address_otherWordsOddChannels_reg <= copy_first_line_others + ROWS_FOR_TILE*row_copy_to + KERNEL*ROWS_FOR_TILE*counter_internal_phase_7 + counter_internal_phase_8 - 3;
            write_address_otherWordsEvenChannels_reg <= copy_first_line_others + ROWS_FOR_TILE*row_copy_to + KERNEL*ROWS_FOR_TILE*counter_internal_phase_7 + counter_internal_phase_8 - 3;
            write_address_firstWordsOddChannels_reg <= copy_first_line_first_six + row_copy_to + KERNEL*counter_internal_phase_7;
            write_address_firstWordsEvenChannels_reg <= copy_first_line_first_six + row_copy_to + KERNEL*counter_internal_phase_7;
            end
        else 
            begin
                if (counter_internal_phase_7 != 0)
                    begin
                    write_address_otherWordsOddChannels_reg <= copy_first_line_others + ROWS_FOR_TILE*row_copy_to + KERNEL*ROWS_FOR_TILE*(counter_internal_phase_7-1) + counter_internal_phase_8 + 4;
                    write_address_otherWordsEvenChannels_reg <= copy_first_line_others + ROWS_FOR_TILE*row_copy_to + KERNEL*ROWS_FOR_TILE*(counter_internal_phase_7-1) + counter_internal_phase_8 + 4;
                    end
            end
    end   
    if (start10 == 1)
        begin
        write_otherWordsEvenChannels_reg <= 0;
        start_copy_row <= 1;
        start10 <= 0;
        start11 <= 1;
        copy_amount_of_channels <= 4;
        copy_first_line_others <= 0;
        copy_first_line_first_six <= 0;
        row_copy_from <= 6;
        row_copy_to <= 0;
        end
    if (start11 == 1)
        if (start_copy_row == 0)
            begin
            start_copy_row <= 1;
            start11 <= 0;
            start12 <= 1;
            copy_amount_of_channels <= 4;
            copy_first_line_others <= 0;
            copy_first_line_first_six <= 0;
            row_copy_from <= 5;
            row_copy_to <= 1;
            end
    if (start12 == 1)
        if (start_copy_row == 0)
            begin
            start_copy_row <= 1;
            start12 <= 0;
            start13 <= 1;
            copy_amount_of_channels <= 4;
            copy_first_line_others <= 0;
            copy_first_line_first_six <= 0;
            row_copy_from <= 4;
            row_copy_to <= 2;
            end
    if (start13 == 1)
        begin
        if (start_copy_row == 0)
            begin
            startFSM <= 1;
            start13 <= 0;
            end
        end
    if (startFSM == 1)
        begin
        case(counterFSM)
        0   :   begin
                startUseful <= 1;
                pointer <= 0;
                first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 3;
                first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 3);
                layer <= 0;
                counterFSM <= counterFSM + 1;
                end
        1   :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        2   :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 1;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 4;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 4);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        3   :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        4   :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 2;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 5;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 5);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        5   :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        6   :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 3;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 6;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 6);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        7   :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER1;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*HALF_CHANNELS_LAYER0;
                    copy_first_line_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    row_copy_from <= 6;
                    row_copy_to <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        8   :   begin
                if (start_copy_row == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER1;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*HALF_CHANNELS_LAYER0;
                    copy_first_line_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    row_copy_from <= 5;
                    row_copy_to <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        9   :   begin
                if (start_copy_row == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER1;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*HALF_CHANNELS_LAYER0;
                    copy_first_line_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    row_copy_from <= 4;
                    row_copy_to <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        10  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 0;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3);
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        11  :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        12  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 4;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        13  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 1;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4);
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        14  :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        15  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 5;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 1;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 1);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        16  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 2;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5);
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        17  :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        18  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 6;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 2;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 2);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        19  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 3;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6);
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        20  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER2;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    row_copy_from <= 6;
                    row_copy_to <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        21  :   begin
                if (start_copy_row == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER2;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    row_copy_from <= 5;
                    row_copy_to <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        22  :   begin
                if (start_copy_row == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER2;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    row_copy_from <= 4;
                    row_copy_to <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        23  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 0;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        24  :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        25  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 0;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 3;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 3);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        26  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 4;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1));
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        27  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 1;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        28  :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        29  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 1;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 4;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 4);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        30  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 5;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1);
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        31  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 2;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        32  :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        33  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 2;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 5;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 5);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        34  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 6;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2);
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        35  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 3;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        36  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER3;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    row_copy_from <= 6;
                    row_copy_to <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        37  :   begin
                if (start_copy_row == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER3;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    row_copy_from <= 5;
                    row_copy_to <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        38  :   begin
                if (start_copy_row == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER3;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    row_copy_from <= 4;
                    row_copy_to <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        39  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 0;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        40  :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        41  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 3;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 6;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 6);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        42  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 0;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3);
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        43  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 4;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        44  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 1;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        45  :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        46  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 4;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        47  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 1;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4);
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        48  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 5;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        49  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 2;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        50  :   begin
                if (startUseful == 0)
                    begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        51  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 5;
                    first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 1;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 1);
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        52  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 2;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5);
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        53  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 6;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        54  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 3;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        55  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER4;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    row_copy_from <= 6;
                    row_copy_to <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        56  :   begin
                if (start_copy_row == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER4;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    row_copy_from <= 5;
                    row_copy_to <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        57  :   begin
                if (start_copy_row == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER4;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    row_copy_from <= 4;
                    row_copy_to <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        58  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    pointer <= 0;
                    first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    pointer1 <= 5;
                    pointer2 <= 2;
                    pointer3 <= 6;
                    pointer4 <= 3;
                    pointer5 <= 0;
                    end
                end
        59  :   begin
                    start_read_new_row <= 1;
                    counterFSM <= counterFSM + 1;
                end
        60  :   begin
                if (start_read_new_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer1 == 6)
                        begin
                        pointer <= 0;
                        pointer1 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer1 + 1;
                        pointer1 <= pointer1 + 1;
                        end
                    case(pointer1)
                    0   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 4;
                    1   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 5;
                    2   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 6;
                    3   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    4   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 1;
                    5   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 2;
                    6   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 3;
                    endcase
                    case(pointer1)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0);
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 3);
                    endcase
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        61  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer2 == 6)
                        begin
                        pointer <= 0;
                        pointer2 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer2 + 1;
                        pointer2 <= pointer2 + 1;
                        end
                    case(pointer2)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3;
                    endcase
                    case(pointer2)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3);
                    endcase
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        62  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        63  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        64  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    case(last_row)
                    0   :   counterFSM <= 59;
                    1   :   counterFSM <= counterFSM + 1;
                    endcase//l
                    end
                end
        65  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER0;
                    copy_first_line_others <= 0;
                    copy_first_line_first_six <= 0;
                    if (pointer1 < 2)
                        row_copy_from <= pointer1 + 5;
                    else
                        row_copy_from <= pointer1 - 2;
                    row_copy_to <= pointer1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        66  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer1 == 6)
                        begin
                        pointer <= 0;
                        pointer1 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer1 + 1;
                        pointer1 <= pointer1 + 1;
                        end
                    case(pointer1)
                    0   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 4;
                    1   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 5;
                    2   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 6;
                    3   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    4   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 1;
                    5   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 2;
                    6   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 3;
                    endcase
                    case(pointer1)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0);
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 3);
                    endcase
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        67  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer2 == 6)
                        begin
                        pointer <= 0;
                        pointer2 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer2 + 1;
                        pointer2 <= pointer2 + 1;
                        end
                    case(pointer2)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3;
                    endcase
                    case(pointer2)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3);
                    endcase
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        68  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        69  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        70  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        71  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER0;
                    copy_first_line_others <= 0;
                    copy_first_line_first_six <= 0;
                    if (pointer1 < 4)
                        row_copy_from <= pointer1 + 3;
                    else
                        row_copy_from <= pointer1 - 4;
                    row_copy_to <= pointer1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        72  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer1 == 6)
                        begin
                        pointer <= 0;
                        pointer1 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer1 + 1;
                        pointer1 <= pointer1 + 1;
                        end
                    case(pointer1)
                    0   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 4;
                    1   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 5;
                    2   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 6;
                    3   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    4   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 1;
                    5   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 2;
                    6   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 3;
                    endcase
                    case(pointer1)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0);
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 3);
                    endcase
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        73  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer2 == 6)
                        begin
                        pointer <= 0;
                        pointer2 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer2 + 1;
                        pointer2 <= pointer2 + 1;
                        end
                    case(pointer2)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3;
                    endcase
                    case(pointer2)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3);
                    endcase
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        74  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        75  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        76  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        77  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER0;
                    copy_first_line_others <= 0;
                    copy_first_line_first_six <= 0;
                    if (pointer1 < 6)
                        row_copy_from <= pointer1 + 1;
                    else
                        row_copy_from <= pointer1 - 6;
                    row_copy_to <= pointer1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        78  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer1 == 6)
                        begin
                        pointer <= 0;
                        pointer1 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer1 + 1;
                        pointer1 <= pointer1 + 1;
                        end
                    case(pointer1)
                    0   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 4;
                    1   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 5;
                    2   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 6;
                    3   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    4   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 1;
                    5   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 2;
                    6   :   first_row_writing_first_six <= KERNEL*HALF_CHANNELS_LAYER0 + 3;
                    endcase
                    case(pointer1)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0);
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*HALF_CHANNELS_LAYER0 + 3);
                    endcase
                    layer <= 0;
                    counterFSM <= counterFSM + 1;
                    end
                end
        79  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer2 == 6)
                        begin
                        pointer <= 0;
                        pointer2 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer2 + 1;
                        pointer2 <= pointer2 + 1;
                        end
                    case(pointer2)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3;
                    endcase
                    case(pointer2)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3);
                    endcase
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        80  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        81  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        82  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        83  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER1;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*HALF_CHANNELS_LAYER0;
                    copy_first_line_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    if (pointer2 < 2)
                        row_copy_from <= pointer2 + 5;
                    else
                        row_copy_from <= pointer2 - 2;
                    row_copy_to <= pointer2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        84  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer2 == 6)
                        begin
                        pointer <= 0;
                        pointer2 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer2 + 1;
                        pointer2 <= pointer2 + 1;
                        end
                    case(pointer2)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3;
                    endcase
                    case(pointer2)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3);
                    endcase
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        85  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        86  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        87  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        88  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER1;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*HALF_CHANNELS_LAYER0;
                    copy_first_line_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    if (pointer2 < 4)
                        row_copy_from <= pointer2 + 3;
                    else
                        row_copy_from <= pointer2 - 4;
                    row_copy_to <= pointer2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        89  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer2 == 6)
                        begin
                        pointer <= 0;
                        pointer2 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer2 + 1;
                        pointer2 <= pointer2 + 1;
                        end
                    case(pointer2)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3;
                    endcase
                    case(pointer2)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3);
                    endcase
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        90  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        91  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        92  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        93  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER1;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*HALF_CHANNELS_LAYER0;
                    copy_first_line_first_six <= KERNEL*HALF_CHANNELS_LAYER0;
                    if (pointer2 < 6)
                        row_copy_from <= pointer2 + 1;
                    else
                        row_copy_from <= pointer2 - 6;
                    row_copy_to <= pointer2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        94  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer2 == 6)
                        begin
                        pointer <= 0;
                        pointer2 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer2 + 1;
                        pointer2 <= pointer2 + 1;
                        end
                    case(pointer2)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3;
                    endcase
                    case(pointer2)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + 3);
                    endcase
                    layer <= 1;
                    counterFSM <= counterFSM + 1;
                    end
                end
        95  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        96  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        97  :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        98  :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER2;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    if (pointer3 < 2)
                        row_copy_from <= pointer3 + 5;
                    else
                        row_copy_from <= pointer3 - 1;
                    row_copy_to <= pointer3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        99  :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        100 :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        101 :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        102 :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER2;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    if (pointer3 < 4)
                        row_copy_from <= pointer3 + 3;
                    else
                        row_copy_from <= pointer3 - 4;
                    row_copy_to <= pointer3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        103 :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        104 :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        105 :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        106 :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER2;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                    if (pointer3 < 6)
                        row_copy_from <= pointer3 + 1;
                    else
                        row_copy_from <= pointer3 - 6;
                    row_copy_to <= pointer3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        107 :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer3 == 6)
                        begin
                        pointer <= 0;
                        pointer3 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer3 + 1;
                        pointer3 <= pointer3 + 1;
                        end
                    case(pointer3)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3;
                    endcase
                    case(pointer3)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + 3);
                    endcase
                    layer <= 2;
                    counterFSM <= counterFSM + 1;
                    end
                end
        108 :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        109 :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        110 :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER3;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    if (pointer4 < 2)
                        row_copy_from <= pointer4 + 5;
                    else
                        row_copy_from <= pointer4 - 2;
                    row_copy_to <= pointer4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        111 :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        112 :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        113 :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER3;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    if (pointer4 < 4)
                        row_copy_from <= pointer4 + 3;
                    else
                        row_copy_from <= pointer4 - 4;
                    row_copy_to <= pointer4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        114 :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        115 :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        116 :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER3;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                    if (pointer4 < 6)
                        row_copy_from <= pointer4 + 1;
                    else
                        row_copy_from <= pointer4 - 6;
                    row_copy_to <= pointer4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        117 :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer4 == 6)
                        begin
                        pointer <= 0;
                        pointer4 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer4 + 1;
                        pointer4 <= pointer4 + 1;
                        end
                    case(pointer4)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3;
                    endcase
                    case(pointer4)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + 3);
                    endcase
                    layer <= 3;
                    counterFSM <= counterFSM + 1;
                    end
                end
        118 :   begin
                if (startUseful == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        119 :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER4;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    if (pointer5 < 2)
                        row_copy_from <= pointer5 + 5;
                    else
                        row_copy_from <= pointer5 - 2;
                    row_copy_to <= pointer5;
                    counterFSM <= counterFSM + 1;
                    end
                end
        120 :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        121 :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER4;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    if (pointer5 < 4)
                        row_copy_from <= pointer5 + 3;
                    else
                        row_copy_from <= pointer5 - 4;
                    row_copy_to <= pointer5;
                    counterFSM <= counterFSM + 1;
                    end
                end
        122 :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        123 :   begin
                if (startUseful == 0)
                    begin
                    start_copy_row <= 1;
                    copy_amount_of_channels <= HALF_CHANNELS_LAYER4;
                    copy_first_line_others <= ROWS_FOR_TILE*KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    copy_first_line_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                    if (pointer5 < 6)
                        row_copy_from <= pointer5 + 1;
                    else
                        row_copy_from <= pointer5 - 6;
                    row_copy_to <= pointer5;
                    counterFSM <= counterFSM + 1;
                    end
                end
        124 :   begin
                if (start_copy_row == 0)
                    begin
                    startUseful <= 1;
                    if (pointer5 == 6)
                        begin
                        pointer <= 0;
                        pointer5 <= 0;
                        end
                    else
                        begin
                        pointer <= pointer5 + 1;
                        pointer5 <= pointer5 + 1;
                        end
                    case(pointer5)
                    0   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4;
                    1   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5;
                    2   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6;
                    3   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4);
                    4   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1;
                    5   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2;
                    6   :   first_row_writing_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3;
                    endcase
                    case(pointer5)
                    0   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 4);
                    1   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 5);
                    2   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 6);
                    3   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4));
                    4   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 1);
                    5   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 2);
                    6   :   first_row_writing_others <= ROWS_FOR_TILE*(KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3+HALF_CHANNELS_LAYER4) + 3);
                    endcase
                    layer <= 4;
                    counterFSM <= counterFSM + 1;
                    end
                end
        125 :   begin
                if (startUseful == 0)
                    done_reg <= 1;
                end
        endcase
        end
    
    // START IMPORTANT
    if (startUseful == 1'b1)
        begin
            case(counter_first_phase)       
            0 : begin  
                counter_internal_phase <= 0;
                counter_internal_phase_1 <= 0;
                counter_internal_phase_2 <= 0;
                counter_internal_phase_3 <= 0;
                case(layer)
                0   :   begin
                        shift_bias <= shift_bias_layer0;  
                        shift_result <= shift_result_layer0;
                        first_row_data_first_six <= 0;
                        first_row_data_others <= 0;
                        first_row_weights <= 0;
                        first_row_biases <= 0;
                        read_address_biasesMemory_reg <= 0; 
                        read_address_weightsOddInputChannelOddOutputChannel_reg <= 0;  
                        read_address_weightsOddInputChannelEvenOutputChannel_reg <= 0;  
                        read_address_weightsEvenInputChannelOddOutputChannel_reg <= 0;  
                        read_address_weightsEvenInputChannelEvenOutputChannel_reg <= 0;   
                        read_address_firstWordsOddChannels_reg <= pointer;
                        read_address_firstWordsEvenChannels_reg <= pointer;
                        number_two_inputs <= HALF_CHANNELS_LAYER0;
                        number_two_outputs <= HALF_CHANNELS_LAYER1;
                        end
                1   :   begin
                        shift_bias <= shift_bias_layer1;  
                        shift_result <= shift_result_layer1;
                        first_row_data_first_six <= KERNEL*(HALF_CHANNELS_LAYER0);
                        first_row_data_others <= KERNEL*ROWS_FOR_TILE*(HALF_CHANNELS_LAYER0);
                        first_row_weights <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1);
                        first_row_biases <= HALF_CHANNELS_LAYER1;
                        read_address_biasesMemory_reg <= HALF_CHANNELS_LAYER1; 
                        read_address_weightsOddInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1);  
                        read_address_weightsOddInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1);  
                        read_address_weightsEvenInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1);  
                        read_address_weightsEvenInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1);   
                        read_address_firstWordsOddChannels_reg <= KERNEL*(HALF_CHANNELS_LAYER0) + pointer;
                        read_address_firstWordsEvenChannels_reg <= KERNEL*(HALF_CHANNELS_LAYER0) + pointer;
                        number_two_inputs <= HALF_CHANNELS_LAYER1;
                        number_two_outputs <= HALF_CHANNELS_LAYER2;
                        end
                2   :   begin
                        shift_bias <= shift_bias_layer2;  
                        shift_result <= shift_result_layer2;
                        first_row_data_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                        first_row_data_others <= KERNEL*ROWS_FOR_TILE*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1);
                        first_row_weights <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2);
                        first_row_biases <= HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER2;
                        read_address_biasesMemory_reg <= HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER2; 
                        read_address_weightsOddInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2);  
                        read_address_weightsOddInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2);  
                        read_address_weightsEvenInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2);  
                        read_address_weightsEvenInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2);   
                        read_address_firstWordsOddChannels_reg <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + pointer;
                        read_address_firstWordsEvenChannels_reg <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1) + pointer;
                        number_two_inputs <= HALF_CHANNELS_LAYER2;
                        number_two_outputs <= HALF_CHANNELS_LAYER3;
                        end
                3   :   begin
                        shift_bias <= shift_bias_layer3;  
                        shift_result <= shift_result_layer3;
                        first_row_data_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                        first_row_data_others <= KERNEL*ROWS_FOR_TILE*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2);
                        first_row_weights <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3);
                        first_row_biases <= HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER3;
                        read_address_biasesMemory_reg <= HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER3; 
                        read_address_weightsOddInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3);  
                        read_address_weightsOddInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3);  
                        read_address_weightsEvenInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3);  
                        read_address_weightsEvenInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3);   
                        read_address_firstWordsOddChannels_reg <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + pointer;
                        read_address_firstWordsEvenChannels_reg <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2) + pointer;
                        number_two_inputs <= HALF_CHANNELS_LAYER3;
                        number_two_outputs <= HALF_CHANNELS_LAYER4;
                        end
                4   :   begin
                        shift_bias <= shift_bias_layer4;  
                        shift_result <= shift_result_layer4;
                        first_row_data_first_six <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                        first_row_data_others <= KERNEL*ROWS_FOR_TILE*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3);
                        first_row_weights <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 
                                                + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4);
                        first_row_biases <= HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER4;
                        read_address_biasesMemory_reg <= HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER3 + HALF_CHANNELS_LAYER4; 
                        read_address_weightsOddInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 
                                                                        + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4);  
                        read_address_weightsOddInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 
                                                                        + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4);  
                        read_address_weightsEvenInputChannelOddOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 
                                                                        + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4);  
                        read_address_weightsEvenInputChannelEvenOutputChannel_reg <= KERNEL*(HALF_CHANNELS_LAYER0*HALF_CHANNELS_LAYER1 + HALF_CHANNELS_LAYER1*HALF_CHANNELS_LAYER2 + HALF_CHANNELS_LAYER2*HALF_CHANNELS_LAYER3 
                                                                        + HALF_CHANNELS_LAYER3*HALF_CHANNELS_LAYER4);   
                        read_address_firstWordsOddChannels_reg <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + pointer;
                        read_address_firstWordsEvenChannels_reg <= KERNEL*(HALF_CHANNELS_LAYER0+HALF_CHANNELS_LAYER1+HALF_CHANNELS_LAYER2+HALF_CHANNELS_LAYER3) + pointer;
                        number_two_inputs <= HALF_CHANNELS_LAYER4;
                        number_two_outputs <= HALF_CHANNELS_LAYER5;
                        end
                endcase
                counter_first_phase <= 1;
                end
            1 : begin
                if (shift_bias == 0)
                    begin
                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer;
                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer;
                    end
                counter_first_phase <= 2;
                end
            2 : begin
                if (shift_bias == 0)
                    begin
                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 1;
                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 1;
                    end
                else if (shift_bias == 1)
                    begin
                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer;
                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer;
                    end
                counter_first_phase <= 3;
                end
            3 : begin
                if (shift_bias == 0)
                    begin
                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 2;
                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 2;
                    end
                else if (shift_bias == 1)
                    begin
                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 1;
                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 1;
                    end
                else if (shift_bias == 2)
                    begin
                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer;
                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer;
                    end
                counter_first_phase <= 4;
                filter_weights_reg <= {weightsOddInputChannelOddOutputChannel_output[KERNEL*BITS-1:0],
                                        weightsEvenInputChannelOddOutputChannel_output[KERNEL*BITS-1:0],
                                        weightsOddInputChannelOddOutputChannel_output[KERNEL*BITS-1:0],
                                        weightsEvenInputChannelOddOutputChannel_output[KERNEL*BITS-1:0],
                                        weightsOddInputChannelEvenOutputChannel_output[KERNEL*BITS-1:0],
                                        weightsEvenInputChannelEvenOutputChannel_output[KERNEL*BITS-1:0],
                                        weightsOddInputChannelEvenOutputChannel_output[KERNEL*BITS-1:0],
                                        weightsEvenInputChannelEvenOutputChannel_output[KERNEL*BITS-1:0]};
                bias_temp1 <= {{(BITS+OVERHEAD_BITS){biasesMemory_output[2*BITS-1]}},biasesMemory_output[2*BITS-1:BITS]};
                bias_temp2 <= {{(BITS+OVERHEAD_BITS){biasesMemory_output[BITS-1]}},biasesMemory_output[BITS-1:0]};
                counter_internal_phase_9 <= 0;
                end
            4 : begin
                if (counter_internal_phase_9 == shift_bias)
                    begin
                    counter_first_phase <= 5;
                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 3;
                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 3;
                    temp_in_1 <= {firstWordsOddChannels_output[(KERNEL-1)*BITS-1:0],otherWordsOddChannels_output[2*(FEATURES-KERNEL+1)*BITS-1:0]};
                    temp_in_2 <= {firstWordsEvenChannels_output[(KERNEL-1)*BITS-1:0],otherWordsEvenChannels_output[2*(FEATURES-KERNEL+1)*BITS-1:0]};
                    end
                else
                    begin
                    case(shift_bias)
                    1   :   begin
                            read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 2;
                            read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 2;
                            end
                    2   :   begin
                            case(counter_internal_phase_9)
                            0   :   begin
                                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 1;
                                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 1;
                                    end
                            1   :   begin
                                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 2;
                                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 2;
                                    end
                            endcase
                            end
                    endcase
                    if (shift_bias >= 3)
                        begin
                        if (counter_internal_phase_9 == shift_bias - 1)
                            begin
                            read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 2;
                            read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 2;
                            end
                        else if (counter_internal_phase_9 == shift_bias - 2)
                            begin
                            read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + 1;
                            read_address_otherWordsEvenChannels_reg <= first_row_data_others + 7*pointer + 1;
                            end
                        else if (counter_internal_phase_9 == shift_bias - 3)
                            begin
                            read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer;
                            read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer;
                            end
                        end
                    counter_internal_phase_9 <= counter_internal_phase_9 + 1;
                    case(bias_temp1[2*BITS+OVERHEAD_BITS-1])
                    0   :   begin
                            if (bias_temp1[2*BITS+OVERHEAD_BITS-2] == 1)
                                bias_temp1[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                            else
                                bias_temp1[2*BITS+OVERHEAD_BITS-2:0] <= {bias_temp1[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                            end
                    1   :   begin
                            if (bias_temp1[2*BITS+OVERHEAD_BITS-2] == 0)
                                bias_temp1[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                            else
                                bias_temp1[2*BITS+OVERHEAD_BITS-2:0] <= {bias_temp1[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                            end
                    endcase
                    case(bias_temp2[2*BITS+OVERHEAD_BITS-1])
                    0   :   begin
                            if (bias_temp2[2*BITS+OVERHEAD_BITS-2] == 1)
                                bias_temp2[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                            else
                                bias_temp2[2*BITS+OVERHEAD_BITS-2:0] <= {bias_temp2[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                            end
                    1   :   begin
                            if (bias_temp2[2*BITS+OVERHEAD_BITS-2] == 0)
                                bias_temp2[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                            else
                                bias_temp2[2*BITS+OVERHEAD_BITS-2:0] <= {bias_temp2[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                            end
                    endcase
                    end
                end
            5 : begin
                if (counter_internal_phase == 0)
                    if (counter_internal_phase_1 == KERNEL - 1)
                        begin
                        if (counter_internal_phase_2 == number_two_inputs - 1)
                            begin
                            read_address_weightsOddInputChannelOddOutputChannel_reg <= first_row_weights + KERNEL*(counter_internal_phase_3 + 1)*number_two_inputs;
                            read_address_weightsOddInputChannelEvenOutputChannel_reg <= first_row_weights + KERNEL*(counter_internal_phase_3 + 1)*number_two_inputs;
                            read_address_weightsEvenInputChannelOddOutputChannel_reg <= first_row_weights + KERNEL*(counter_internal_phase_3 + 1)*number_two_inputs;
                            read_address_weightsEvenInputChannelEvenOutputChannel_reg <= first_row_weights + KERNEL*(counter_internal_phase_3 + 1)*number_two_inputs;
                            end    
                        else
                            begin
                            read_address_weightsOddInputChannelOddOutputChannel_reg <= first_row_weights + KERNEL*counter_internal_phase_3*number_two_inputs + KERNEL*counter_internal_phase_2 + 1 + counter_internal_phase_1;
                            read_address_weightsOddInputChannelEvenOutputChannel_reg <= first_row_weights + KERNEL*counter_internal_phase_3*number_two_inputs + KERNEL*counter_internal_phase_2 + 1 + counter_internal_phase_1;
                            read_address_weightsEvenInputChannelOddOutputChannel_reg <= first_row_weights + KERNEL*counter_internal_phase_3*number_two_inputs + KERNEL*counter_internal_phase_2 + 1 + counter_internal_phase_1;
                            read_address_weightsEvenInputChannelEvenOutputChannel_reg <= first_row_weights + KERNEL*counter_internal_phase_3*number_two_inputs + KERNEL*counter_internal_phase_2 + 1 + counter_internal_phase_1;
                            end    
                        end
                    else
                        begin
                        read_address_weightsOddInputChannelOddOutputChannel_reg <= first_row_weights + KERNEL*counter_internal_phase_3*number_two_inputs + KERNEL*counter_internal_phase_2 + 1 + counter_internal_phase_1;
                        read_address_weightsOddInputChannelEvenOutputChannel_reg <= first_row_weights + KERNEL*counter_internal_phase_3*number_two_inputs + KERNEL*counter_internal_phase_2 + 1 + counter_internal_phase_1;
                        read_address_weightsEvenInputChannelOddOutputChannel_reg <= first_row_weights + KERNEL*counter_internal_phase_3*number_two_inputs + KERNEL*counter_internal_phase_2 + 1 + counter_internal_phase_1;
                        read_address_weightsEvenInputChannelEvenOutputChannel_reg <= first_row_weights + KERNEL*counter_internal_phase_3*number_two_inputs + KERNEL*counter_internal_phase_2 + 1 + counter_internal_phase_1;
                        end
                if (counter_internal_phase_2 == 0)
                    begin
                        if (counter_internal_phase_1 == 0)
                            begin
                            biases_reg[54*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:53*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1){bias_temp1}};
                            biases_reg[47*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:46*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                            biases_reg[36*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:35*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1){bias_temp1}};
                            biases_reg[35*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:34*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                            biases_reg[26*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:25*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1){bias_temp2}};
                            biases_reg[19*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:18*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                            biases_reg[8*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:7*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1){bias_temp2}};
                            biases_reg[7*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:6*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                            if (counter_internal_phase == 5)
                                begin
                                    biases_reg_temp_2 <= results;
                                end
                            if (counter_internal_phase == 6)
                                begin
                                    biases_reg_temp_2 <= results;
                                    biases_reg_temp_1 <= biases_reg_temp_2;
                                end
                            end
                        else
                            begin
                                biases_reg[54*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:53*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= biases_reg_temp_1[4*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:3*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)];
                                biases_reg[47*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:46*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                                biases_reg[36*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:35*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= biases_reg_temp_1[3*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:2*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)];
                                biases_reg[35*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:34*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                                biases_reg[26*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:25*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= biases_reg_temp_1[2*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)];
                                biases_reg[19*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:18*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                                biases_reg[8*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:7*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= biases_reg_temp_1[(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0];
                                biases_reg[7*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:6*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                                biases_reg_temp_1 <= biases_reg_temp_2;
                                biases_reg_temp_2 <= results;
                            end
                    end
                else
                    begin
                    read_address_biasesMemory_reg <= first_row_biases + counter_internal_phase_3 + 1;
                    biases_reg[54*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:53*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= biases_reg_temp_1[4*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:3*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)];
                    biases_reg[47*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:46*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                    biases_reg[36*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:35*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= biases_reg_temp_1[3*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:2*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)];
                    biases_reg[35*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:34*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                    biases_reg[26*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:25*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= biases_reg_temp_1[2*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)];
                    biases_reg[19*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:18*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                    biases_reg[8*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:7*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= biases_reg_temp_1[(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:0];
                    biases_reg[7*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)-1:6*(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS)] <= {(FEATURES-KERNEL+1)*(2*BITS+OVERHEAD_BITS){1'b0}};
                    biases_reg_temp_1 <= biases_reg_temp_2;
                    biases_reg_temp_2 <= results;
                    end
                if (counter_internal_phase_2 == 1)
                    if (counter_internal_phase_1 == 0)
                        if (counter_internal_phase == 3)
                            begin
                            bias_temp1 <= {{(BITS+OVERHEAD_BITS){biasesMemory_output[2*BITS-1]}},biasesMemory_output[2*BITS-1:BITS]};
                            bias_temp2 <= {{(BITS+OVERHEAD_BITS){biasesMemory_output[BITS-1]}},biasesMemory_output[BITS-1:0]};
                            counter_internal_phase_9 <= 0;
                            end
                if (counter_internal_phase_9 != shift_bias)
                    begin
                    counter_internal_phase_9 <= counter_internal_phase_9 + 1;
                    case(bias_temp1[2*BITS+OVERHEAD_BITS-1])
                    0   :   begin
                            if (bias_temp1[2*BITS+OVERHEAD_BITS-2] == 1)
                                bias_temp1[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                            else
                                bias_temp1[2*BITS+OVERHEAD_BITS-2:0] <= {bias_temp1[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                            end
                    1   :   begin
                            if (bias_temp1[2*BITS+OVERHEAD_BITS-2] == 0)
                                bias_temp1[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                            else
                                bias_temp1[2*BITS+OVERHEAD_BITS-2:0] <= {bias_temp1[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                            end
                    endcase
                    case(bias_temp2[2*BITS+OVERHEAD_BITS-1])
                    0   :   begin
                            if (bias_temp2[2*BITS+OVERHEAD_BITS-2] == 1)
                                bias_temp2[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                            else
                                bias_temp2[2*BITS+OVERHEAD_BITS-2:0] <= {bias_temp2[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                            end
                    1   :   begin
                            if (bias_temp2[2*BITS+OVERHEAD_BITS-2] == 0)
                                bias_temp2[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                            else
                                bias_temp2[2*BITS+OVERHEAD_BITS-2:0] <= {bias_temp2[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                            end
                    endcase
                    end
                if (counter_internal_phase < 3)
                    begin
                        if (pointer + counter_internal_phase_1 >= KERNEL)
                            begin
                                read_address_otherWordsOddChannels_reg <= first_row_data_others + KERNEL*ROWS_FOR_TILE*counter_internal_phase_2 + ROWS_FOR_TILE*(pointer + counter_internal_phase_1 - KERNEL) + counter_internal_phase + 4;
                                read_address_otherWordsEvenChannels_reg <= first_row_data_others + KERNEL*ROWS_FOR_TILE*counter_internal_phase_2 + ROWS_FOR_TILE*(pointer + counter_internal_phase_1 - KERNEL) + counter_internal_phase + 4;
                            end
                        else
                            begin
                                read_address_otherWordsOddChannels_reg <= first_row_data_others + KERNEL*ROWS_FOR_TILE*counter_internal_phase_2 + ROWS_FOR_TILE*(pointer + counter_internal_phase_1) + counter_internal_phase + 4;
                                read_address_otherWordsEvenChannels_reg <= first_row_data_others + KERNEL*ROWS_FOR_TILE*counter_internal_phase_2 + ROWS_FOR_TILE*(pointer + counter_internal_phase_1) + counter_internal_phase + 4;
                            end
                    end  
                else
                    begin
                        if (counter_internal_phase_1 == KERNEL - 1)
                            begin
                                if (counter_internal_phase_2 == number_two_inputs - 1)
                                    begin
                                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + counter_internal_phase - 3;
                                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*pointer + counter_internal_phase - 3;
                                    end
                                else
                                    begin
                                    read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*KERNEL*(counter_internal_phase_2+1) + ROWS_FOR_TILE*pointer + counter_internal_phase - 3;
                                    read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*KERNEL*(counter_internal_phase_2+1) + ROWS_FOR_TILE*pointer + counter_internal_phase - 3;
                                    end
                            end
                        else
                            begin
                                if (pointer + counter_internal_phase_1 + 1 >= KERNEL)
                                    begin
                                        read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*KERNEL*counter_internal_phase_2 + ROWS_FOR_TILE*(pointer + counter_internal_phase_1 - KERNEL + 1) + counter_internal_phase - 3;
                                        read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*KERNEL*counter_internal_phase_2 + ROWS_FOR_TILE*(pointer + counter_internal_phase_1 - KERNEL + 1) + counter_internal_phase - 3;
                                    end
                                else
                                    begin
                                        read_address_otherWordsOddChannels_reg <= first_row_data_others + ROWS_FOR_TILE*KERNEL*counter_internal_phase_2 + ROWS_FOR_TILE*(pointer + counter_internal_phase_1 + 1) + counter_internal_phase - 3;
                                        read_address_otherWordsEvenChannels_reg <= first_row_data_others + ROWS_FOR_TILE*KERNEL*counter_internal_phase_2 + ROWS_FOR_TILE*(pointer + counter_internal_phase_1 + 1) + counter_internal_phase - 3;
                                    end
                            end
                    end
                if (counter_internal_phase == 3)
                    begin
                        if (counter_internal_phase_1 == KERNEL - 1)
                            begin
                                if (counter_internal_phase_2 == number_two_inputs - 1)
                                    begin
                                    read_address_firstWordsOddChannels_reg <= first_row_data_first_six + pointer;
                                    read_address_firstWordsEvenChannels_reg <= first_row_data_first_six + pointer;
                                    end
                                else
                                    begin
                                    read_address_firstWordsOddChannels_reg <= first_row_data_first_six + pointer + KERNEL*(counter_internal_phase_2+1);
                                    read_address_firstWordsEvenChannels_reg <= first_row_data_first_six + pointer + KERNEL*(counter_internal_phase_2+1);
                                    end
                            end
                        else
                            begin
                                if (pointer + counter_internal_phase_1 + 1 >= KERNEL)
                                    begin
                                        read_address_firstWordsOddChannels_reg <= first_row_data_first_six + (pointer+counter_internal_phase_1-KERNEL+1) + KERNEL*counter_internal_phase_2;
                                        read_address_firstWordsEvenChannels_reg <= first_row_data_first_six + (pointer+counter_internal_phase_1-KERNEL+1) + KERNEL*counter_internal_phase_2;
                                    end
                                else
                                    begin
                                        read_address_firstWordsOddChannels_reg <= first_row_data_first_six + (pointer+counter_internal_phase_1+1) + KERNEL*counter_internal_phase_2;
                                        read_address_firstWordsEvenChannels_reg <= first_row_data_first_six + (pointer+counter_internal_phase_1+1) + KERNEL*counter_internal_phase_2;
                                    end
                            end
                    end                                       
                if (counter_internal_phase == ROWS_FOR_TILE - 1)
                    begin
                    temp_in_1 <= {firstWordsOddChannels_output[(KERNEL-1)*BITS-1:0],otherWordsOddChannels_output[2*(FEATURES-KERNEL+1)*BITS-1:0]};
                    temp_in_2 <= {firstWordsEvenChannels_output[(KERNEL-1)*BITS-1:0],otherWordsEvenChannels_output[2*(FEATURES-KERNEL+1)*BITS-1:0]};
                    end
                else
                    begin
                    temp_in_1 <= {temp_in_1[(KERNEL-1)*BITS-1:0],otherWordsOddChannels_output[2*(FEATURES-KERNEL+1)*BITS-1:0]};
                    temp_in_2 <= {temp_in_2[(KERNEL-1)*BITS-1:0],otherWordsEvenChannels_output[2*(FEATURES-KERNEL+1)*BITS-1:0]};
                    end                          
                if (counter_internal_phase == ROWS_FOR_TILE - 1)
                    begin
                        filter_weights_reg <= {weightsOddInputChannelOddOutputChannel_output[KERNEL*BITS-1:0],
                                                weightsEvenInputChannelOddOutputChannel_output[KERNEL*BITS-1:0],
                                                weightsOddInputChannelOddOutputChannel_output[KERNEL*BITS-1:0],
                                                weightsEvenInputChannelOddOutputChannel_output[KERNEL*BITS-1:0],
                                                weightsOddInputChannelEvenOutputChannel_output[KERNEL*BITS-1:0],
                                                weightsEvenInputChannelEvenOutputChannel_output[KERNEL*BITS-1:0],
                                                weightsOddInputChannelEvenOutputChannel_output[KERNEL*BITS-1:0],
                                                weightsEvenInputChannelEvenOutputChannel_output[KERNEL*BITS-1:0]};
                        counter_internal_phase <= 0;
                        if (counter_internal_phase_1 == KERNEL - 1)
                            begin
                                counter_internal_phase_1 <= 0;
                                if (counter_internal_phase_2 == number_two_inputs - 1)
                                    begin
                                        counter_internal_phase_2 <= 0;
                                        if (counter_internal_phase_3 == number_two_outputs - 1)
                                            begin
                                            counter_internal_phase_3 <= 0;
                                            counter_first_phase <= 6;
                                            end
                                        else
                                            counter_internal_phase_3 <= counter_internal_phase_3 + 1;
                                    end
                                else
                                    counter_internal_phase_2 <= counter_internal_phase_2 + 1;
                            end
                        else
                            counter_internal_phase_1 <= counter_internal_phase_1 + 1;
                    end//for
                else
                    counter_internal_phase <= counter_internal_phase + 1;
                if (counter_internal_phase_2 == number_two_inputs - 1)
                    if (counter_internal_phase_1 == KERNEL - 1)
                        if (counter_internal_phase == 4)
                            counter_internal_phase_4 <= 0;
                end
            6 : begin
                if (counter_internal_phase_4 == 16)
                    begin
                    startUseful <= 0;
                    counter_first_phase <= 0;
                    end
                end
            endcase
  end
  
  // END IMPORTANT
  case(counter_internal_phase_4)   
  0  :  begin
        if (type[2] == 1)
            begin
                results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-1:174*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-1:0] <= {(174*(2*BITS+OVERHEAD_BITS)){1'b0}};
                results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-1:174*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
                results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-1:0] <= {(174*(2*BITS+OVERHEAD_BITS)){1'b0}};
            end
        else
            begin
                results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-1:203*(2*BITS+OVERHEAD_BITS)] <= results[57*(2*BITS+OVERHEAD_BITS)-1:56*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-1:202*(2*BITS+OVERHEAD_BITS)] <= results[58*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-1:201*(2*BITS+OVERHEAD_BITS)] <= results[59*(2*BITS+OVERHEAD_BITS)-1:58*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-1:171*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-1:0] <= {(171*(2*BITS+OVERHEAD_BITS)){1'b0}};
                results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-1:203*(2*BITS+OVERHEAD_BITS)] <= results[27*(2*BITS+OVERHEAD_BITS)-1:26*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-1:202*(2*BITS+OVERHEAD_BITS)] <= results[28*(2*BITS+OVERHEAD_BITS)-1:27*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-1:201*(2*BITS+OVERHEAD_BITS)] <= results[29*(2*BITS+OVERHEAD_BITS)-1:28*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-1:171*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
                results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-1:0] <= {(171*(2*BITS+OVERHEAD_BITS)){1'b0}};
            end
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
  1 :   begin
        if (type[2] == 1)
            begin
                results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-1:144*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-1:144*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
            end
        else
            begin
                results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-1:141*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-1:141*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
            end
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
  2  :  begin
        if (type[2] == 1)
            begin
                results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-1:114*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-1:114*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
            end
        else
            begin
                results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-1:111*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-1:111*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
            end
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
    3 : begin
        if (type[2] == 1)
            begin
                results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-1:84*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-1:84*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
            end
        else
            begin
                results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-1:81*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-1:81*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
            end
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
    4 : begin
        if (type[2] == 1)
            begin
                results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
            end
        else
            begin
                results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
            end
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
    5 : begin
            if (type[2] == 1)
                begin
                    results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                    results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:0];
                    if (type == 6)
                        begin
                        if (layer == 4)
                            begin
                            results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-1:23*(2*BITS+OVERHEAD_BITS)] <= results[32*(2*BITS+OVERHEAD_BITS)-1:31*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-1:22*(2*BITS+OVERHEAD_BITS)] <= results[33*(2*BITS+OVERHEAD_BITS)-1:32*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)] <= results[34*(2*BITS+OVERHEAD_BITS)-1:33*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-1:23*(2*BITS+OVERHEAD_BITS)] <= results[2*(2*BITS+OVERHEAD_BITS)-1:(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-1:22*(2*BITS+OVERHEAD_BITS)] <= results[3*(2*BITS+OVERHEAD_BITS)-1:2*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)] <= results[4*(2*BITS+OVERHEAD_BITS)-1:3*(2*BITS+OVERHEAD_BITS)];
                            end
                        else if (layer == 3)
                            begin
                            results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[31*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[(2*BITS+OVERHEAD_BITS)-1:0];
                            end
                        end
                end
            else
                begin
                    results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-1:41*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:50*(2*BITS+OVERHEAD_BITS)];
                    results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-1:41*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)];
                    if (type == 0)
                        begin
                        results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-1:40*(2*BITS+OVERHEAD_BITS)] <= results[52*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)];
                        results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-1:39*(2*BITS+OVERHEAD_BITS)] <= results[53*(2*BITS+OVERHEAD_BITS)-1:52*(2*BITS+OVERHEAD_BITS)];
                        results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-1:38*(2*BITS+OVERHEAD_BITS)] <= results[54*(2*BITS+OVERHEAD_BITS)-1:53*(2*BITS+OVERHEAD_BITS)];
                        results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-1:40*(2*BITS+OVERHEAD_BITS)] <= results[22*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)];
                        results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-1:39*(2*BITS+OVERHEAD_BITS)] <= results[23*(2*BITS+OVERHEAD_BITS)-1:22*(2*BITS+OVERHEAD_BITS)];
                        results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-1:38*(2*BITS+OVERHEAD_BITS)] <= results[24*(2*BITS+OVERHEAD_BITS)-1:23*(2*BITS+OVERHEAD_BITS)];
                        end
                    else
                        begin
                            results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)] <= results[50*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)] <= results[20*(2*BITS+OVERHEAD_BITS)-1:0];
                            if (type == 1)
                                begin
                                results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)] <= results[32*(2*BITS+OVERHEAD_BITS)-1:31*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-1:19*(2*BITS+OVERHEAD_BITS)] <= results[33*(2*BITS+OVERHEAD_BITS)-1:32*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[34*(2*BITS+OVERHEAD_BITS)-1:33*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)] <= results[2*(2*BITS+OVERHEAD_BITS)-1:(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-1:19*(2*BITS+OVERHEAD_BITS)] <= results[3*(2*BITS+OVERHEAD_BITS)-1:2*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[4*(2*BITS+OVERHEAD_BITS)-1:3*(2*BITS+OVERHEAD_BITS)];
                                end
                        end
                end
            counter_internal_phase_4 <= counter_internal_phase_4 + 1;
            end
    6  :    begin
            case(type)
            2   :   begin
                    if (layer != 4)
                        begin
                        results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)];
                        results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:27*(2*BITS+OVERHEAD_BITS)];
                        if (layer != 3)
                            begin
                            results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-1:15*(2*BITS+OVERHEAD_BITS)] <= results[57*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-1:15*(2*BITS+OVERHEAD_BITS)] <= results[27*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)];
                            if (layer != 2)
                                begin
                                results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)] <= results[54*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)] <= results[24*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)];
                                if (layer == 0)
                                    begin
                                    results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-1:9*(2*BITS+OVERHEAD_BITS)] <= results[51*(2*BITS+OVERHEAD_BITS)-1:48*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-1:9*(2*BITS+OVERHEAD_BITS)] <= results[21*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)];
                                    end
                                end
                            end
                        end
                    end
            4   :   begin
                    if (layer != 4)
                        begin
                        results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)];
                        results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)];
                        if (layer != 3)
                            begin
                            results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)] <= results[54*(2*BITS+OVERHEAD_BITS)-1:48*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)] <= results[24*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)];
                            if (layer != 2)
                                begin
                                results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-1:6*(2*BITS+OVERHEAD_BITS)] <= results[48*(2*BITS+OVERHEAD_BITS)-1:42*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-1:6*(2*BITS+OVERHEAD_BITS)] <= results[18*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)];
                                if (layer == 0)
                                    begin
                                    results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-1:0] <= results[42*(2*BITS+OVERHEAD_BITS)-1:36*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-1:0] <= results[12*(2*BITS+OVERHEAD_BITS)-1:6*(2*BITS+OVERHEAD_BITS)];
                                    end
                                end
                            end
                        end
                    end
            6   :   begin
                    if (layer != 4)
                        begin
                        results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)];
                        results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:27*(2*BITS+OVERHEAD_BITS)];
                        if (layer != 3)
                            begin
                            results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[57*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)] <= results[27*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)];
                            if (layer != 2)
                                begin
                                results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-1:15*(2*BITS+OVERHEAD_BITS)] <= results[54*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-1:15*(2*BITS+OVERHEAD_BITS)] <= results[24*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)];
                                if (layer == 0)
                                    begin
                                    results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)] <= results[51*(2*BITS+OVERHEAD_BITS)-1:48*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)] <= results[21*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-1:11*(2*BITS+OVERHEAD_BITS)] <= results[50*(2*BITS+OVERHEAD_BITS)-1:49*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-1:10*(2*BITS+OVERHEAD_BITS)] <= results[51*(2*BITS+OVERHEAD_BITS)-1:50*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-1:9*(2*BITS+OVERHEAD_BITS)] <= results[52*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-1:11*(2*BITS+OVERHEAD_BITS)] <= results[20*(2*BITS+OVERHEAD_BITS)-1:19*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-1:10*(2*BITS+OVERHEAD_BITS)] <= results[21*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-1:9*(2*BITS+OVERHEAD_BITS)] <= results[22*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)];
                                    end
                                else
                                    begin
                                    results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-1:14*(2*BITS+OVERHEAD_BITS)] <= results[53*(2*BITS+OVERHEAD_BITS)-1:52*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-1:13*(2*BITS+OVERHEAD_BITS)] <= results[54*(2*BITS+OVERHEAD_BITS)-1:53*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)] <= results[55*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-1:14*(2*BITS+OVERHEAD_BITS)] <= results[23*(2*BITS+OVERHEAD_BITS)-1:22*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-1:13*(2*BITS+OVERHEAD_BITS)] <= results[24*(2*BITS+OVERHEAD_BITS)-1:23*(2*BITS+OVERHEAD_BITS)];
                                    results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)] <= results[25*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)];
                                    end
                                end
                            else
                                begin
                                results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-1:17*(2*BITS+OVERHEAD_BITS)] <= results[56*(2*BITS+OVERHEAD_BITS)-1:55*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-1:16*(2*BITS+OVERHEAD_BITS)] <= results[57*(2*BITS+OVERHEAD_BITS)-1:56*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-1:15*(2*BITS+OVERHEAD_BITS)] <= results[58*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-1:17*(2*BITS+OVERHEAD_BITS)] <= results[26*(2*BITS+OVERHEAD_BITS)-1:25*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-1:16*(2*BITS+OVERHEAD_BITS)] <= results[27*(2*BITS+OVERHEAD_BITS)-1:26*(2*BITS+OVERHEAD_BITS)];
                                results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-1:15*(2*BITS+OVERHEAD_BITS)] <= results[28*(2*BITS+OVERHEAD_BITS)-1:27*(2*BITS+OVERHEAD_BITS)];
                                end
                            end
                        else
                            begin
                            results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)] <= results[59*(2*BITS+OVERHEAD_BITS)-1:58*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-1:19*(2*BITS+OVERHEAD_BITS)] <= results[60*(2*BITS+OVERHEAD_BITS)-1:59*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)] <= results[29*(2*BITS+OVERHEAD_BITS)-1:28*(2*BITS+OVERHEAD_BITS)];
                            results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-1:19*(2*BITS+OVERHEAD_BITS)] <= results[30*(2*BITS+OVERHEAD_BITS)-1:29*(2*BITS+OVERHEAD_BITS)];
                            end
                        end
                    end
            endcase
            counter_internal_phase_4 <= counter_internal_phase_4 + 1;
            counter_internal_phase_10 <= 0;
        end
  7 :   begin
        if (counter_internal_phase_10 != shift_result)
            begin
            counter_internal_phase_10 <= counter_internal_phase_10 + 1;
            case(results_to_write_in_ram_1[2*BITS+OVERHEAD_BITS-1])
            0   :   case(results_to_write_in_ram_1[2*BITS+OVERHEAD_BITS-2])
                    1   :   results_to_write_in_ram_1[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[2*BITS+OVERHEAD_BITS-2:0] <= {results_to_write_in_ram_1[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[2*BITS+OVERHEAD_BITS-2])
                    0   :   results_to_write_in_ram_1[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[2*BITS+OVERHEAD_BITS-2:0] <= {results_to_write_in_ram_1[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-2:2*BITS+OVERHEAD_BITS] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-2:2*BITS+OVERHEAD_BITS] <= {results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-3:2*BITS+OVERHEAD_BITS],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-2:2*BITS+OVERHEAD_BITS] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-2:2*BITS+OVERHEAD_BITS] <= {results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-3:2*BITS+OVERHEAD_BITS],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-2:2*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-2:2*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-3:2*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-2:2*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-2:2*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-3:2*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-2:3*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-2:3*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-3:3*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-2:3*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-2:3*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-3:3*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-2:4*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-2:4*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-3:4*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-2:4*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-2:4*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-3:4*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-2:5*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-2:5*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-3:5*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-2:5*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-2:5*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-3:5*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-2:6*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-2:6*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-3:6*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-2:6*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-2:6*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-3:6*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-2:7*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-2:7*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-3:7*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-2:7*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-2:7*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-3:7*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-2:8*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-2:8*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-3:8*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-2:8*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-2:8*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-3:8*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-2:9*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-2:9*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-3:9*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-2:9*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-2:9*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-3:9*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-2:10*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-2:10*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-3:10*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-2:10*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-2:10*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-3:10*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-2:11*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-2:11*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-3:11*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-2:11*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-2:11*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-3:11*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-2:12*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-2:12*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-3:12*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-2:12*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-2:12*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-3:12*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-2:13*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-2:13*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-3:13*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-2:13*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-2:13*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-3:13*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-2:14*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-2:14*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-3:14*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-2:14*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-2:14*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-3:14*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-2:15*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-2:15*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-3:15*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-2:15*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-2:15*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-3:15*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-2:16*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-2:16*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-3:16*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-2:16*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-2:16*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-3:16*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-2:17*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-2:17*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-3:17*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-2:17*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-2:17*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-3:17*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-2:18*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-2:18*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-3:18*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-2:18*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-2:18*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-3:18*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-2:19*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-2:19*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-3:19*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-2:19*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-2:19*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-3:19*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-2:20*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-2:20*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-3:20*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-2:20*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-2:20*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-3:20*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-2:21*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-2:21*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-3:21*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-2:21*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-2:21*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-3:21*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-2:22*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-2:22*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-3:22*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-2:22*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-2:22*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-3:22*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-2:23*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-2:23*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-3:23*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-2:23*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-2:23*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-3:23*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-2:24*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-2:24*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-3:24*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-2:24*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-2:24*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-3:24*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-2:25*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-2:25*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-3:25*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-2:25*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-2:25*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-3:25*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-2:26*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-2:26*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-3:26*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-2:26*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-2:26*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-3:26*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-2:27*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-2:27*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-3:27*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-2:27*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-2:27*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-3:27*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-2:28*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-2:28*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-3:28*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-2:28*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-2:28*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-3:28*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-2:29*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-2:29*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-3:29*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-2:29*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-2:29*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-3:29*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-2:30*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-2:30*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-3:30*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-2:30*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-2:30*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-3:30*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-2:31*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-2:31*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-3:31*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-2:31*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-2:31*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-3:31*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-2:32*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-2:32*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-3:32*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-2:32*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-2:32*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-3:32*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-2:33*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-2:33*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-3:33*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-2:33*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-2:33*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-3:33*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-2:34*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-2:34*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-3:34*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-2:34*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-2:34*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-3:34*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-2:35*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-2:35*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-3:35*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-2:35*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-2:35*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-3:35*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-2:36*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-2:36*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-3:36*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-2:36*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-2:36*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-3:36*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-2:37*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-2:37*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-3:37*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-2:37*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-2:37*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-3:37*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-2:38*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-2:38*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-3:38*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-2:38*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-2:38*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-3:38*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-2:39*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-2:39*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-3:39*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-2:39*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-2:39*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-3:39*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-2:40*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-2:40*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-3:40*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-2:40*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-2:40*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-3:40*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-2:41*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-2:41*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-3:41*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-2:41*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-2:41*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-3:41*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-2:42*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-2:42*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-3:42*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-2:42*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-2:42*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-3:42*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-2:43*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-2:43*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-3:43*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-2:43*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-2:43*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-3:43*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-2:44*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-2:44*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-3:44*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-2:44*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-2:44*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-3:44*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-2:45*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-2:45*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-3:45*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-2:45*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-2:45*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-3:45*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-2:46*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-2:46*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-3:46*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-2:46*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-2:46*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-3:46*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-2:47*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-2:47*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-3:47*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-2:47*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-2:47*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-3:47*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-2:48*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-2:48*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-3:48*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-2:48*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-2:48*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-3:48*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-2:49*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-2:49*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-3:49*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-2:49*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-2:49*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-3:49*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-2:50*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-2:50*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-3:50*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-2:50*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-2:50*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-3:50*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-2:51*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-2:51*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-3:51*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-2:51*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-2:51*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-3:51*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-2:52*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-2:52*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-3:52*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-2:52*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-2:52*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-3:52*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-2:53*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-2:53*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-3:53*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-2:53*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-2:53*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-3:53*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-2:54*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-2:54*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-3:54*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-2:54*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-2:54*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-3:54*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-2:55*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-2:55*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-3:55*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-2:55*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-2:55*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-3:55*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-2:56*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-2:56*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-3:56*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-2:56*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-2:56*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-3:56*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-2:57*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-2:57*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-3:57*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-2:57*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-2:57*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-3:57*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-2:58*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-2:58*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-3:58*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-2:58*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-2:58*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-3:58*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-2:59*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-2:59*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-3:59*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-2:59*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-2:59*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-3:59*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-2:60*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-2:60*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-3:60*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-2:60*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-2:60*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-3:60*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-2:61*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-2:61*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-3:61*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-2:61*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-2:61*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-3:61*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-2:62*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-2:62*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-3:62*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-2:62*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-2:62*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-3:62*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-2:63*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-2:63*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-3:63*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-2:63*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-2:63*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-3:63*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-2:64*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-2:64*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-3:64*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-2:64*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-2:64*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-3:64*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-2:65*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-2:65*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-3:65*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-2:65*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-2:65*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-3:65*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-2:66*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-2:66*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-3:66*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-2:66*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-2:66*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-3:66*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-2:67*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-2:67*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-3:67*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-2:67*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-2:67*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-3:67*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-2:68*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-2:68*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-3:68*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-2:68*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-2:68*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-3:68*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-2:69*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-2:69*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-3:69*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-2:69*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-2:69*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-3:69*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-2:70*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-2:70*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-3:70*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-2:70*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-2:70*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-3:70*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-2:71*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-2:71*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-3:71*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-2:71*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-2:71*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-3:71*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-2:72*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-2:72*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-3:72*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-2:72*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-2:72*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-3:72*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-2:73*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-2:73*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-3:73*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-2:73*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-2:73*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-3:73*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-2:74*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-2:74*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-3:74*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-2:74*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-2:74*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-3:74*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-2:75*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-2:75*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-3:75*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-2:75*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-2:75*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-3:75*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-2:76*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-2:76*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-3:76*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-2:76*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-2:76*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-3:76*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-2:77*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-2:77*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-3:77*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-2:77*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-2:77*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-3:77*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-2:78*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-2:78*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-3:78*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-2:78*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-2:78*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-3:78*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-2:79*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-2:79*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-3:79*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-2:79*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-2:79*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-3:79*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-2:80*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-2:80*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-3:80*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-2:80*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-2:80*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-3:80*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-2:81*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-2:81*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-3:81*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-2:81*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-2:81*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-3:81*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-2:82*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-2:82*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-3:82*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-2:82*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-2:82*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-3:82*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-2:83*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-2:83*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-3:83*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-2:83*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-2:83*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-3:83*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-2:84*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-2:84*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-3:84*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-2:84*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-2:84*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-3:84*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-2:85*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-2:85*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-3:85*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-2:85*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-2:85*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-3:85*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-2:86*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-2:86*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-3:86*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-2:86*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-2:86*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-3:86*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-2:87*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-2:87*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-3:87*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-2:87*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-2:87*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-3:87*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-2:88*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-2:88*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-3:88*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-2:88*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-2:88*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-3:88*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-2:89*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-2:89*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-3:89*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-2:89*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-2:89*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-3:89*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-2:90*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-2:90*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-3:90*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-2:90*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-2:90*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-3:90*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-2:91*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-2:91*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-3:91*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-2:91*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-2:91*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-3:91*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-2:92*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-2:92*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-3:92*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-2:92*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-2:92*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-3:92*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-2:93*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-2:93*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-3:93*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-2:93*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-2:93*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-3:93*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-2:94*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-2:94*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-3:94*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-2:94*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-2:94*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-3:94*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-2:95*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-2:95*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-3:95*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-2:95*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-2:95*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-3:95*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-2:96*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-2:96*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-3:96*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-2:96*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-2:96*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-3:96*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-2:97*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-2:97*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-3:97*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-2:97*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-2:97*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-3:97*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-2:98*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-2:98*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-3:98*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-2:98*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-2:98*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-3:98*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-2:99*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-2:99*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-3:99*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-2:99*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-2:99*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-3:99*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-2:100*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-2:100*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-3:100*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-2:100*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-2:100*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-3:100*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-2:101*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-2:101*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-3:101*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-2:101*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-2:101*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-3:101*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-2:102*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-2:102*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-3:102*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-2:102*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-2:102*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-3:102*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-2:103*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-2:103*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-3:103*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-2:103*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-2:103*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-3:103*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-2:104*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-2:104*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-3:104*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-2:104*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-2:104*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-3:104*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-2:105*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-2:105*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-3:105*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-2:105*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-2:105*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-3:105*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-2:106*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-2:106*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-3:106*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-2:106*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-2:106*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-3:106*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-2:107*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-2:107*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-3:107*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-2:107*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-2:107*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-3:107*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-2:108*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-2:108*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-3:108*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-2:108*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-2:108*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-3:108*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-2:109*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-2:109*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-3:109*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-2:109*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-2:109*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-3:109*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-2:110*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-2:110*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-3:110*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-2:110*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-2:110*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-3:110*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-2:111*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-2:111*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-3:111*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-2:111*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-2:111*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-3:111*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-2:112*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-2:112*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-3:112*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-2:112*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-2:112*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-3:112*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-2:113*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-2:113*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-3:113*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-2:113*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-2:113*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-3:113*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-2:114*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-2:114*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-3:114*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-2:114*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-2:114*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-3:114*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-2:115*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-2:115*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-3:115*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-2:115*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-2:115*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-3:115*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-2:116*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-2:116*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-3:116*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-2:116*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-2:116*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-3:116*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-2:117*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-2:117*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-3:117*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-2:117*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-2:117*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-3:117*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-2:118*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-2:118*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-3:118*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-2:118*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-2:118*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-3:118*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-2:119*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-2:119*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-3:119*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-2:119*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-2:119*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-3:119*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-2:120*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-2:120*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-3:120*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-2:120*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-2:120*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-3:120*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-2:121*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-2:121*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-3:121*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-2:121*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-2:121*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-3:121*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-2:122*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-2:122*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-3:122*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-2:122*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-2:122*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-3:122*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-2:123*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-2:123*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-3:123*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-2:123*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-2:123*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-3:123*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-2:124*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-2:124*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-3:124*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-2:124*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-2:124*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-3:124*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-2:125*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-2:125*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-3:125*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-2:125*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-2:125*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-3:125*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-2:126*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-2:126*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-3:126*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-2:126*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-2:126*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-3:126*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-2:127*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-2:127*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-3:127*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-2:127*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-2:127*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-3:127*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-2:128*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-2:128*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-3:128*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-2:128*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-2:128*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-3:128*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-2:129*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-2:129*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-3:129*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-2:129*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-2:129*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-3:129*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-2:130*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-2:130*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-3:130*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-2:130*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-2:130*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-3:130*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-2:131*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-2:131*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-3:131*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-2:131*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-2:131*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-3:131*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-2:132*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-2:132*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-3:132*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-2:132*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-2:132*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-3:132*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-2:133*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-2:133*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-3:133*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-2:133*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-2:133*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-3:133*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-2:134*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-2:134*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-3:134*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-2:134*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-2:134*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-3:134*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-2:135*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-2:135*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-3:135*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-2:135*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-2:135*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-3:135*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-2:136*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-2:136*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-3:136*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-2:136*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-2:136*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-3:136*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-2:137*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-2:137*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-3:137*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-2:137*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-2:137*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-3:137*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-2:138*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-2:138*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-3:138*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-2:138*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-2:138*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-3:138*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-2:139*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-2:139*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-3:139*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-2:139*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-2:139*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-3:139*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-2:140*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-2:140*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-3:140*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-2:140*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-2:140*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-3:140*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-2:141*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-2:141*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-3:141*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-2:141*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-2:141*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-3:141*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-2:142*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-2:142*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-3:142*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-2:142*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-2:142*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-3:142*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-2:143*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-2:143*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-3:143*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-2:143*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-2:143*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-3:143*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-2:144*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-2:144*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-3:144*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-2:144*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-2:144*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-3:144*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-2:145*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-2:145*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-3:145*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-2:145*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-2:145*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-3:145*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-2:146*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-2:146*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-3:146*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-2:146*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-2:146*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-3:146*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-2:147*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-2:147*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-3:147*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-2:147*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-2:147*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-3:147*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-2:148*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-2:148*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-3:148*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-2:148*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-2:148*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-3:148*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-2:149*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-2:149*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-3:149*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-2:149*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-2:149*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-3:149*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-2:150*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-2:150*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-3:150*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-2:150*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-2:150*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-3:150*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-2:151*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-2:151*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-3:151*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-2:151*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-2:151*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-3:151*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-2:152*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-2:152*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-3:152*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-2:152*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-2:152*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-3:152*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-2:153*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-2:153*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-3:153*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-2:153*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-2:153*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-3:153*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-2:154*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-2:154*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-3:154*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-2:154*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-2:154*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-3:154*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-2:155*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-2:155*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-3:155*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-2:155*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-2:155*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-3:155*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-2:156*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-2:156*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-3:156*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-2:156*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-2:156*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-3:156*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-2:157*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-2:157*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-3:157*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-2:157*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-2:157*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-3:157*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-2:158*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-2:158*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-3:158*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-2:158*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-2:158*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-3:158*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-2:159*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-2:159*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-3:159*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-2:159*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-2:159*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-3:159*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-2:160*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-2:160*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-3:160*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-2:160*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-2:160*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-3:160*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-2:161*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-2:161*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-3:161*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-2:161*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-2:161*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-3:161*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-2:162*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-2:162*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-3:162*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-2:162*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-2:162*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-3:162*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-2:163*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-2:163*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-3:163*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-2:163*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-2:163*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-3:163*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-2:164*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-2:164*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-3:164*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-2:164*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-2:164*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-3:164*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-2:165*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-2:165*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-3:165*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-2:165*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-2:165*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-3:165*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-2:166*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-2:166*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-3:166*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-2:166*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-2:166*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-3:166*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-2:167*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-2:167*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-3:167*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-2:167*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-2:167*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-3:167*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-2:168*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-2:168*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-3:168*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-2:168*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-2:168*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-3:168*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-2:169*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-2:169*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-3:169*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-2:169*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-2:169*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-3:169*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-2:170*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-2:170*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-3:170*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-2:170*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-2:170*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-3:170*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-2:171*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-2:171*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-3:171*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-2:171*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-2:171*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-3:171*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-2:172*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-2:172*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-3:172*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-2:172*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-2:172*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-3:172*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-2:173*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-2:173*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-3:173*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-2:173*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-2:173*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-3:173*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-2:174*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-2:174*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-3:174*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-2:174*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-2:174*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-3:174*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-2:175*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-2:175*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-3:175*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-2:175*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-2:175*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-3:175*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-2:176*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-2:176*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-3:176*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-2:176*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-2:176*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-3:176*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-2:177*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-2:177*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-3:177*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-2:177*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-2:177*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-3:177*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-2:178*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-2:178*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-3:178*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-2:178*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-2:178*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-3:178*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-2:179*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-2:179*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-3:179*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-2:179*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-2:179*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-3:179*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-2:180*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-2:180*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-3:180*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-2:180*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-2:180*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-3:180*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-2:181*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-2:181*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-3:181*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-2:181*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-2:181*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-3:181*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-2:182*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-2:182*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-3:182*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-2:182*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-2:182*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-3:182*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-2:183*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-2:183*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-3:183*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-2:183*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-2:183*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-3:183*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-2:184*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-2:184*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-3:184*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-2:184*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-2:184*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-3:184*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-2:185*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-2:185*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-3:185*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-2:185*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-2:185*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-3:185*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-2:186*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-2:186*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-3:186*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-2:186*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-2:186*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-3:186*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-2:187*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-2:187*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-3:187*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-2:187*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-2:187*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-3:187*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-2:188*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-2:188*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-3:188*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-2:188*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-2:188*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-3:188*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-2:189*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-2:189*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-3:189*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-2:189*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-2:189*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-3:189*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-2:190*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-2:190*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-3:190*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-2:190*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-2:190*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-3:190*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-2:191*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-2:191*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-3:191*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-2:191*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-2:191*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-3:191*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-2:192*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-2:192*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-3:192*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-2:192*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-2:192*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-3:192*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-2:193*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-2:193*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-3:193*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-2:193*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-2:193*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-3:193*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-2:194*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-2:194*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-3:194*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-2:194*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-2:194*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-3:194*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-2:195*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-2:195*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-3:195*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-2:195*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-2:195*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-3:195*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-2:196*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-2:196*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-3:196*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-2:196*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-2:196*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-3:196*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-2:197*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-2:197*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-3:197*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-2:197*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-2:197*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-3:197*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-2:198*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-2:198*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-3:198*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-2:198*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-2:198*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-3:198*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-2:199*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-2:199*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-3:199*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-2:199*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-2:199*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-3:199*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-2:200*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-2:200*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-3:200*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-2:200*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-2:200*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-3:200*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-2:201*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-2:201*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-3:201*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-2:201*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-2:201*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-3:201*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-2:202*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-2:202*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-3:202*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-2:202*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-2:202*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-3:202*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-2:203*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-2:203*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-3:203*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-2:203*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-2:203*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-3:203*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[2*BITS+OVERHEAD_BITS-1])
            0   :   case(results_to_write_in_ram_2[2*BITS+OVERHEAD_BITS-2])
                    1   :   results_to_write_in_ram_2[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[2*BITS+OVERHEAD_BITS-2:0] <= {results_to_write_in_ram_2[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[2*BITS+OVERHEAD_BITS-2])
                    0   :   results_to_write_in_ram_2[2*BITS+OVERHEAD_BITS-2:0] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[2*BITS+OVERHEAD_BITS-2:0] <= {results_to_write_in_ram_2[2*BITS+OVERHEAD_BITS-3:0],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-2:2*BITS+OVERHEAD_BITS] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-2:2*BITS+OVERHEAD_BITS] <= {results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-3:2*BITS+OVERHEAD_BITS],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-2:2*BITS+OVERHEAD_BITS] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-2:2*BITS+OVERHEAD_BITS] <= {results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-3:2*BITS+OVERHEAD_BITS],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-2:2*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-2:2*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-3:2*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-2:2*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-2:2*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-3:2*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-2:3*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-2:3*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-3:3*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-2:3*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-2:3*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-3:3*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-2:4*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-2:4*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-3:4*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-2:4*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-2:4*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-3:4*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-2:5*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-2:5*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-3:5*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-2:5*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-2:5*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-3:5*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-2:6*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-2:6*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-3:6*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-2:6*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-2:6*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-3:6*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-2:7*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-2:7*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-3:7*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-2:7*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-2:7*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-3:7*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-2:8*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-2:8*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-3:8*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-2:8*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-2:8*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-3:8*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-2:9*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-2:9*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-3:9*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-2:9*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-2:9*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-3:9*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-2:10*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-2:10*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-3:10*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-2:10*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-2:10*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-3:10*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-2:11*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-2:11*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-3:11*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-2:11*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-2:11*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-3:11*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-2:12*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-2:12*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-3:12*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-2:12*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-2:12*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-3:12*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-2:13*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-2:13*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-3:13*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-2:13*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-2:13*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-3:13*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-2:14*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-2:14*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-3:14*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-2:14*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-2:14*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-3:14*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-2:15*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-2:15*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-3:15*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-2:15*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-2:15*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-3:15*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-2:16*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-2:16*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-3:16*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-2:16*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-2:16*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-3:16*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-2:17*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-2:17*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-3:17*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-2:17*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-2:17*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-3:17*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-2:18*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-2:18*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-3:18*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-2:18*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-2:18*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-3:18*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-2:19*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-2:19*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-3:19*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-2:19*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-2:19*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-3:19*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-2:20*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-2:20*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-3:20*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-2:20*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-2:20*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-3:20*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-2:21*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-2:21*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-3:21*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-2:21*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-2:21*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-3:21*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-2:22*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-2:22*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-3:22*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-2:22*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-2:22*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-3:22*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-2:23*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-2:23*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-3:23*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-2:23*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-2:23*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-3:23*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-2:24*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-2:24*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-3:24*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-2:24*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-2:24*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-3:24*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-2:25*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-2:25*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-3:25*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-2:25*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-2:25*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-3:25*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-2:26*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-2:26*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-3:26*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-2:26*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-2:26*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-3:26*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-2:27*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-2:27*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-3:27*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-2:27*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-2:27*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-3:27*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-2:28*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-2:28*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-3:28*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-2:28*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-2:28*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-3:28*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-2:29*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-2:29*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-3:29*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-2:29*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-2:29*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-3:29*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-2:30*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-2:30*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-3:30*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-2:30*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-2:30*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-3:30*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-2:31*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-2:31*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-3:31*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-2:31*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-2:31*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-3:31*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-2:32*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-2:32*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-3:32*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-2:32*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-2:32*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-3:32*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-2:33*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-2:33*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-3:33*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-2:33*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-2:33*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-3:33*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-2:34*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-2:34*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-3:34*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-2:34*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-2:34*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-3:34*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-2:35*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-2:35*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-3:35*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-2:35*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-2:35*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-3:35*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-2:36*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-2:36*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-3:36*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-2:36*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-2:36*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-3:36*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-2:37*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-2:37*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-3:37*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-2:37*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-2:37*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-3:37*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-2:38*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-2:38*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-3:38*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-2:38*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-2:38*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-3:38*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-2:39*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-2:39*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-3:39*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-2:39*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-2:39*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-3:39*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-2:40*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-2:40*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-3:40*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-2:40*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-2:40*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-3:40*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-2:41*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-2:41*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-3:41*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-2:41*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-2:41*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-3:41*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-2:42*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-2:42*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-3:42*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-2:42*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-2:42*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-3:42*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-2:43*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-2:43*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-3:43*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-2:43*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-2:43*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-3:43*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-2:44*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-2:44*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-3:44*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-2:44*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-2:44*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-3:44*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-2:45*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-2:45*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-3:45*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-2:45*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-2:45*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-3:45*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-2:46*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-2:46*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-3:46*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-2:46*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-2:46*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-3:46*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-2:47*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-2:47*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-3:47*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-2:47*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-2:47*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-3:47*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-2:48*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-2:48*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-3:48*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-2:48*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-2:48*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-3:48*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-2:49*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-2:49*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-3:49*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-2:49*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-2:49*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-3:49*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-2:50*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-2:50*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-3:50*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-2:50*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-2:50*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-3:50*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-2:51*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-2:51*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-3:51*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-2:51*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-2:51*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-3:51*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-2:52*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-2:52*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-3:52*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-2:52*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-2:52*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-3:52*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-2:53*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-2:53*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-3:53*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-2:53*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-2:53*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-3:53*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-2:54*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-2:54*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-3:54*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-2:54*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-2:54*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-3:54*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-2:55*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-2:55*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-3:55*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-2:55*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-2:55*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-3:55*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-2:56*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-2:56*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-3:56*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-2:56*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-2:56*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-3:56*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-2:57*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-2:57*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-3:57*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-2:57*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-2:57*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-3:57*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-2:58*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-2:58*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-3:58*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-2:58*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-2:58*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-3:58*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-2:59*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-2:59*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-3:59*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-2:59*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-2:59*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-3:59*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-2:60*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-2:60*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-3:60*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-2:60*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-2:60*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-3:60*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-2:61*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-2:61*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-3:61*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-2:61*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-2:61*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-3:61*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-2:62*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-2:62*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-3:62*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-2:62*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-2:62*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-3:62*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-2:63*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-2:63*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-3:63*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-2:63*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-2:63*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-3:63*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-2:64*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-2:64*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-3:64*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-2:64*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-2:64*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-3:64*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-2:65*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-2:65*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-3:65*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-2:65*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-2:65*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-3:65*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-2:66*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-2:66*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-3:66*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-2:66*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-2:66*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-3:66*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-2:67*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-2:67*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-3:67*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-2:67*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-2:67*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-3:67*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-2:68*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-2:68*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-3:68*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-2:68*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-2:68*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-3:68*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-2:69*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-2:69*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-3:69*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-2:69*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-2:69*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-3:69*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-2:70*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-2:70*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-3:70*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-2:70*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-2:70*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-3:70*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-2:71*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-2:71*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-3:71*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-2:71*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-2:71*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-3:71*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-2:72*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-2:72*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-3:72*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-2:72*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-2:72*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-3:72*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-2:73*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-2:73*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-3:73*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-2:73*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-2:73*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-3:73*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-2:74*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-2:74*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-3:74*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-2:74*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-2:74*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-3:74*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-2:75*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-2:75*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-3:75*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-2:75*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-2:75*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-3:75*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-2:76*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-2:76*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-3:76*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-2:76*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-2:76*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-3:76*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-2:77*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-2:77*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-3:77*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-2:77*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-2:77*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-3:77*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-2:78*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-2:78*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-3:78*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-2:78*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-2:78*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-3:78*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-2:79*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-2:79*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-3:79*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-2:79*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-2:79*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-3:79*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-2:80*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-2:80*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-3:80*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-2:80*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-2:80*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-3:80*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-2:81*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-2:81*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-3:81*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-2:81*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-2:81*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-3:81*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-2:82*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-2:82*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-3:82*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-2:82*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-2:82*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-3:82*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-2:83*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-2:83*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-3:83*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-2:83*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-2:83*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-3:83*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-2:84*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-2:84*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-3:84*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-2:84*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-2:84*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-3:84*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-2:85*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-2:85*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-3:85*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-2:85*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-2:85*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-3:85*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-2:86*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-2:86*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-3:86*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-2:86*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-2:86*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-3:86*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-2:87*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-2:87*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-3:87*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-2:87*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-2:87*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-3:87*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-2:88*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-2:88*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-3:88*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-2:88*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-2:88*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-3:88*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-2:89*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-2:89*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-3:89*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-2:89*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-2:89*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-3:89*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-2:90*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-2:90*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-3:90*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-2:90*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-2:90*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-3:90*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-2:91*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-2:91*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-3:91*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-2:91*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-2:91*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-3:91*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-2:92*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-2:92*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-3:92*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-2:92*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-2:92*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-3:92*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-2:93*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-2:93*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-3:93*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-2:93*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-2:93*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-3:93*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-2:94*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-2:94*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-3:94*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-2:94*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-2:94*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-3:94*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-2:95*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-2:95*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-3:95*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-2:95*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-2:95*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-3:95*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-2:96*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-2:96*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-3:96*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-2:96*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-2:96*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-3:96*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-2:97*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-2:97*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-3:97*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-2:97*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-2:97*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-3:97*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-2:98*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-2:98*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-3:98*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-2:98*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-2:98*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-3:98*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-2:99*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-2:99*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-3:99*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-2:99*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-2:99*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-3:99*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-2:100*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-2:100*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-3:100*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-2:100*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-2:100*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-3:100*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-2:101*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-2:101*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-3:101*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-2:101*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-2:101*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-3:101*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-2:102*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-2:102*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-3:102*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-2:102*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-2:102*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-3:102*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-2:103*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-2:103*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-3:103*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-2:103*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-2:103*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-3:103*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-2:104*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-2:104*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-3:104*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-2:104*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-2:104*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-3:104*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-2:105*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-2:105*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-3:105*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-2:105*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-2:105*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-3:105*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-2:106*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-2:106*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-3:106*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-2:106*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-2:106*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-3:106*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-2:107*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-2:107*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-3:107*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-2:107*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-2:107*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-3:107*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-2:108*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-2:108*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-3:108*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-2:108*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-2:108*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-3:108*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-2:109*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-2:109*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-3:109*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-2:109*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-2:109*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-3:109*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-2:110*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-2:110*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-3:110*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-2:110*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-2:110*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-3:110*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-2:111*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-2:111*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-3:111*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-2:111*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-2:111*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-3:111*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-2:112*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-2:112*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-3:112*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-2:112*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-2:112*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-3:112*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-2:113*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-2:113*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-3:113*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-2:113*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-2:113*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-3:113*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-2:114*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-2:114*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-3:114*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-2:114*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-2:114*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-3:114*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-2:115*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-2:115*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-3:115*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-2:115*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-2:115*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-3:115*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-2:116*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-2:116*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-3:116*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-2:116*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-2:116*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-3:116*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-2:117*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-2:117*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-3:117*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-2:117*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-2:117*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-3:117*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-2:118*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-2:118*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-3:118*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-2:118*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-2:118*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-3:118*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-2:119*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-2:119*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-3:119*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-2:119*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-2:119*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-3:119*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-2:120*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-2:120*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-3:120*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-2:120*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-2:120*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-3:120*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-2:121*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-2:121*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-3:121*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-2:121*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-2:121*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-3:121*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-2:122*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-2:122*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-3:122*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-2:122*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-2:122*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-3:122*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-2:123*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-2:123*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-3:123*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-2:123*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-2:123*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-3:123*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-2:124*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-2:124*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-3:124*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-2:124*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-2:124*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-3:124*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-2:125*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-2:125*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-3:125*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-2:125*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-2:125*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-3:125*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-2:126*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-2:126*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-3:126*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-2:126*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-2:126*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-3:126*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-2:127*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-2:127*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-3:127*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-2:127*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-2:127*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-3:127*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-2:128*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-2:128*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-3:128*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-2:128*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-2:128*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-3:128*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-2:129*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-2:129*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-3:129*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-2:129*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-2:129*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-3:129*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-2:130*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-2:130*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-3:130*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-2:130*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-2:130*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-3:130*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-2:131*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-2:131*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-3:131*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-2:131*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-2:131*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-3:131*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-2:132*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-2:132*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-3:132*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-2:132*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-2:132*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-3:132*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-2:133*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-2:133*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-3:133*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-2:133*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-2:133*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-3:133*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-2:134*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-2:134*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-3:134*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-2:134*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-2:134*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-3:134*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-2:135*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-2:135*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-3:135*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-2:135*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-2:135*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-3:135*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-2:136*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-2:136*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-3:136*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-2:136*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-2:136*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-3:136*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-2:137*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-2:137*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-3:137*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-2:137*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-2:137*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-3:137*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-2:138*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-2:138*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-3:138*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-2:138*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-2:138*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-3:138*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-2:139*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-2:139*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-3:139*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-2:139*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-2:139*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-3:139*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-2:140*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-2:140*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-3:140*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-2:140*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-2:140*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-3:140*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-2:141*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-2:141*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-3:141*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-2:141*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-2:141*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-3:141*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-2:142*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-2:142*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-3:142*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-2:142*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-2:142*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-3:142*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-2:143*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-2:143*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-3:143*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-2:143*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-2:143*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-3:143*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-2:144*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-2:144*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-3:144*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-2:144*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-2:144*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-3:144*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-2:145*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-2:145*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-3:145*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-2:145*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-2:145*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-3:145*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-2:146*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-2:146*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-3:146*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-2:146*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-2:146*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-3:146*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-2:147*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-2:147*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-3:147*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-2:147*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-2:147*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-3:147*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-2:148*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-2:148*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-3:148*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-2:148*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-2:148*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-3:148*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-2:149*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-2:149*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-3:149*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-2:149*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-2:149*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-3:149*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-2:150*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-2:150*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-3:150*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-2:150*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-2:150*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-3:150*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-2:151*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-2:151*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-3:151*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-2:151*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-2:151*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-3:151*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-2:152*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-2:152*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-3:152*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-2:152*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-2:152*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-3:152*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-2:153*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-2:153*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-3:153*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-2:153*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-2:153*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-3:153*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-2:154*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-2:154*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-3:154*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-2:154*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-2:154*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-3:154*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-2:155*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-2:155*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-3:155*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-2:155*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-2:155*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-3:155*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-2:156*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-2:156*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-3:156*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-2:156*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-2:156*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-3:156*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-2:157*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-2:157*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-3:157*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-2:157*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-2:157*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-3:157*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-2:158*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-2:158*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-3:158*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-2:158*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-2:158*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-3:158*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-2:159*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-2:159*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-3:159*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-2:159*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-2:159*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-3:159*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-2:160*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-2:160*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-3:160*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-2:160*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-2:160*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-3:160*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-2:161*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-2:161*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-3:161*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-2:161*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-2:161*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-3:161*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-2:162*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-2:162*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-3:162*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-2:162*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-2:162*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-3:162*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-2:163*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-2:163*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-3:163*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-2:163*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-2:163*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-3:163*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-2:164*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-2:164*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-3:164*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-2:164*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-2:164*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-3:164*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-2:165*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-2:165*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-3:165*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-2:165*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-2:165*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-3:165*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-2:166*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-2:166*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-3:166*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-2:166*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-2:166*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-3:166*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-2:167*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-2:167*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-3:167*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-2:167*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-2:167*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-3:167*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-2:168*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-2:168*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-3:168*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-2:168*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-2:168*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-3:168*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-2:169*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-2:169*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-3:169*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-2:169*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-2:169*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-3:169*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-2:170*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-2:170*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-3:170*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-2:170*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-2:170*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-3:170*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-2:171*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-2:171*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-3:171*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-2:171*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-2:171*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-3:171*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-2:172*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-2:172*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-3:172*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-2:172*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-2:172*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-3:172*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-2:173*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-2:173*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-3:173*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-2:173*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-2:173*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-3:173*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-2:174*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-2:174*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-3:174*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-2:174*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-2:174*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-3:174*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-2:175*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-2:175*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-3:175*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-2:175*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-2:175*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-3:175*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-2:176*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-2:176*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-3:176*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-2:176*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-2:176*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-3:176*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-2:177*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-2:177*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-3:177*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-2:177*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-2:177*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-3:177*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-2:178*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-2:178*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-3:178*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-2:178*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-2:178*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-3:178*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-2:179*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-2:179*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-3:179*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-2:179*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-2:179*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-3:179*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-2:180*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-2:180*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-3:180*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-2:180*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-2:180*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-3:180*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-2:181*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-2:181*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-3:181*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-2:181*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-2:181*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-3:181*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-2:182*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-2:182*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-3:182*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-2:182*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-2:182*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-3:182*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-2:183*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-2:183*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-3:183*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-2:183*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-2:183*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-3:183*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-2:184*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-2:184*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-3:184*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-2:184*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-2:184*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-3:184*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-2:185*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-2:185*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-3:185*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-2:185*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-2:185*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-3:185*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-2:186*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-2:186*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-3:186*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-2:186*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-2:186*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-3:186*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-2:187*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-2:187*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-3:187*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-2:187*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-2:187*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-3:187*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-2:188*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-2:188*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-3:188*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-2:188*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-2:188*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-3:188*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-2:189*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-2:189*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-3:189*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-2:189*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-2:189*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-3:189*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-2:190*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-2:190*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-3:190*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-2:190*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-2:190*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-3:190*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-2:191*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-2:191*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-3:191*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-2:191*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-2:191*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-3:191*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-2:192*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-2:192*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-3:192*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-2:192*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-2:192*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-3:192*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-2:193*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-2:193*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-3:193*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-2:193*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-2:193*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-3:193*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-2:194*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-2:194*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-3:194*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-2:194*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-2:194*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-3:194*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-2:195*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-2:195*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-3:195*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-2:195*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-2:195*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-3:195*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-2:196*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-2:196*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-3:196*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-2:196*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-2:196*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-3:196*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-2:197*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-2:197*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-3:197*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-2:197*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-2:197*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-3:197*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-2:198*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-2:198*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-3:198*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-2:198*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-2:198*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-3:198*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-2:199*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-2:199*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-3:199*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-2:199*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-2:199*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-3:199*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-2:200*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-2:200*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-3:200*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-2:200*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-2:200*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-3:200*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-2:201*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-2:201*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-3:201*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-2:201*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-2:201*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-3:201*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-2:202*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-2:202*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-3:202*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-2:202*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-2:202*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-3:202*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            case(results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-1])
            0   :   case(results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-2])
                    1   :   results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-2:203*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b1}};
                    0   :   results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-2:203*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-3:203*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            1   :   case(results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-2])
                    0   :   results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-2:203*(2*BITS+OVERHEAD_BITS)] <= {(2*BITS+OVERHEAD_BITS-1){1'b0}};
                    1   :   results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-2:203*(2*BITS+OVERHEAD_BITS)] <= {results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-3:203*(2*BITS+OVERHEAD_BITS)],1'b0};
                    endcase
            endcase
            end
        else
            begin
            if (layer != 4)
                counter_internal_phase_4 <= counter_internal_phase_4 + 1;
            else
                begin
                start_to_output <= 1;
                counter_internal_phase_6 <= 0;
                writing_row <= 0;
                end
            end
        end
  8 :   begin
        write_firstWordsOddChannels_reg <= 1;
        write_firstWordsEvenChannels_reg <= 1;
        write_otherWordsOddChannels_reg <= 1;
        write_otherWordsEvenChannels_reg <= 1;
        write_address_firstWordsOddChannels_reg <= first_row_writing_first_six;
        case(results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-1:204*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-1:203*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-1:202*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-1:201*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsOddChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-1:200*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsOddChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsOddChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-1:199*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsOddChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        write_address_firstWordsEvenChannels_reg <= first_row_writing_first_six;
        case(results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-1:204*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-1:203*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-1:202*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-1:201*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsEvenChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-1:200*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsEvenChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-1])
        0   :   firstWordsEvenChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-1:199*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   firstWordsEvenChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        write_address_otherWordsOddChannels_reg <= first_row_writing_others;
        case(results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-1:198*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-1:197*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-1:196*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-1:195*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-1:194*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-1:193*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-1:192*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-1:191*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-1:190*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-1:189*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-1:188*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-1:187*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-1:186*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-1:185*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-1:184*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-1:183*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-1:182*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-1:181*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-1:180*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-1:179*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-1:178*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-1:177*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-1:176*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-1:175*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-1:174*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-1:173*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-1:172*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-1:171*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-1:170*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-1:169*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        write_address_otherWordsEvenChannels_reg <= first_row_writing_others;
        case(results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-1:198*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-1:197*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-1:196*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-1:195*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-1:194*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-1:193*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-1:192*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-1:191*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-1:190*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-1:189*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-1:188*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-1:187*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-1:186*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-1:185*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-1:184*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-1:183*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-1:182*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-1:181*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-1:180*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-1:179*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-1:178*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-1:177*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-1:176*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-1:175*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-1:174*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-1:173*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-1:172*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-1:171*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-1:170*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-1:169*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
  9 :   begin
        write_firstWordsOddChannels_reg <= 0;
        write_firstWordsEvenChannels_reg <= 0;
        first_row_writing_first_six <= first_row_writing_first_six + 7;
        write_address_otherWordsOddChannels_reg <= first_row_writing_others + 1;
        case(results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-1:168*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-1:167*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-1:166*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-1:165*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-1:164*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-1:163*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-1:162*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-1:161*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-1:160*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-1:159*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-1:158*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-1:157*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-1:156*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-1:155*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-1:154*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-1:153*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-1:152*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-1:151*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-1:150*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-1:149*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-1:148*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-1:147*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-1:146*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-1:145*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-1:144*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-1:143*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-1:142*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-1:141*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-1:140*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-1:139*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        write_address_otherWordsEvenChannels_reg <= first_row_writing_others + 1;
        case(results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-1:168*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-1:167*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-1:166*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-1:165*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-1:164*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-1:163*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-1:162*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-1:161*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-1:160*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-1:159*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-1:158*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-1:157*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-1:156*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-1:155*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-1:154*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-1:153*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-1:152*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-1:151*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-1:150*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-1:149*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-1:148*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-1:147*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-1:146*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-1:145*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-1:144*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-1:143*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-1:142*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-1:141*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-1:140*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-1:139*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
  10 :  begin
        write_address_otherWordsOddChannels_reg <= first_row_writing_others + 2;
        case(results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-1:138*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-1:137*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-1:136*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-1:135*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-1:134*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-1:133*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-1:132*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-1:131*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-1:130*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-1:129*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-1:128*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-1:127*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-1:126*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-1:125*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-1:124*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-1:123*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-1:122*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-1:121*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-1:120*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-1:119*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-1:118*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-1:117*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-1:116*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-1:115*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-1:114*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-1:113*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-1:112*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-1:111*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-1:110*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-1:109*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        write_address_otherWordsEvenChannels_reg <= first_row_writing_others + 2;
        case(results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-1:138*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-1:137*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-1:136*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-1:135*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-1:134*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-1:133*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-1:132*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-1:131*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-1:130*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-1:129*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-1:128*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-1:127*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-1:126*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-1:125*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-1:124*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-1:123*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-1:122*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-1:121*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-1:120*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-1:119*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-1:118*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-1:117*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-1:116*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-1:115*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-1:114*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-1:113*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-1:112*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-1:111*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-1:110*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-1:109*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
  11 :  begin
        write_address_otherWordsOddChannels_reg <= first_row_writing_others + 3;
        case(results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-1:108*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-1:107*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-1:106*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-1:105*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-1:104*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-1:103*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-1:102*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-1:101*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-1:100*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-1:99*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-1:98*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-1:97*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-1:96*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-1:95*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-1:94*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-1:93*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-1:92*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-1:91*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-1:90*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-1:89*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-1:88*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-1:87*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-1:86*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-1:85*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-1:84*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-1:83*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-1:82*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-1:81*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-1:80*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-1:79*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        write_address_otherWordsEvenChannels_reg <= first_row_writing_others + 3;
        case(results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-1:108*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-1:107*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-1:106*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-1:105*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-1:104*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-1:103*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-1:102*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-1:101*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-1:100*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-1:99*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-1:98*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-1:97*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-1:96*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-1:95*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-1:94*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-1:93*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-1:92*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-1:91*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-1:90*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-1:89*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-1:88*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-1:87*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-1:86*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-1:85*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-1:84*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-1:83*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-1:82*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-1:81*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-1:80*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-1:79*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
  12 :  begin
        write_address_otherWordsOddChannels_reg <= first_row_writing_others + 4;
        case(results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-1:78*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-1:77*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-1:76*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-1:75*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-1:74*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-1:73*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-1:72*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-1:71*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-1:70*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-1:69*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-1:68*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-1:67*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-1:66*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-1:65*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-1:64*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-1:63*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-1:62*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-1:61*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-1:60*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-1:59*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-1:58*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-1:56*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-1:55*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-1:53*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-1:52*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-1:50*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-1:49*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        write_address_otherWordsEvenChannels_reg <= first_row_writing_others + 4;
        case(results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-1:78*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-1:77*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-1:76*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-1:75*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-1:74*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-1:73*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-1:72*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-1:71*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-1:70*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-1:69*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-1:68*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-1:67*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-1:66*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-1:65*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-1:64*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-1:63*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-1:62*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-1:61*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-1:60*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-1:59*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-1:58*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-1:56*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-1:55*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-1:53*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-1:52*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-1:50*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-1:49*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
  13 :  begin
        write_address_otherWordsOddChannels_reg <= first_row_writing_others + 5;
        case(results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-1:48*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-1:47*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-1:46*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-1:45*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-1:44*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-1:43*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-1:42*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-1:41*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-1:40*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-1:39*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-1:38*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-1:37*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-1:36*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-1:35*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-1:34*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-1:33*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-1:32*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-1:31*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-1:29*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-1:28*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-1:27*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-1:26*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-1:25*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-1:23*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-1:22*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-1:19*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        write_address_otherWordsEvenChannels_reg <= first_row_writing_others + 5;
        case(results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-1:48*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-1:47*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-1:46*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-1:45*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-1:44*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-1:43*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-1:42*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-1:41*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-1:40*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-1:39*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-1:38*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-1:37*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-1:36*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-1:35*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-1:34*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-1:33*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-1:32*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-1:31*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[12*BITS-1:11*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-1:29*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[11*BITS-1:10*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-1:28*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[10*BITS-1:9*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-1:27*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[9*BITS-1:8*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-1:26*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[8*BITS-1:7*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-1:25*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[7*BITS-1:6*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[6*BITS-1:5*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-1:23*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[5*BITS-1:4*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-1:22*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[4*BITS-1:3*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[3*BITS-1:2*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[2*BITS-1:BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-1:19*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[BITS-1:0] <= {BITS{1'b0}};
        endcase
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
  14 :  begin
        write_address_otherWordsOddChannels_reg <= first_row_writing_others + 6;
        case(results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_1[18*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_1[17*(2*BITS+OVERHEAD_BITS)-1:17*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_1[16*(2*BITS+OVERHEAD_BITS)-1:16*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_1[15*(2*BITS+OVERHEAD_BITS)-1:15*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_1[14*(2*BITS+OVERHEAD_BITS)-1:14*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_1[13*(2*BITS+OVERHEAD_BITS)-1:13*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_1[12*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_1[11*(2*BITS+OVERHEAD_BITS)-1:11*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_1[10*(2*BITS+OVERHEAD_BITS)-1:10*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_1[9*(2*BITS+OVERHEAD_BITS)-1:9*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_1[8*(2*BITS+OVERHEAD_BITS)-1:8*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_1[7*(2*BITS+OVERHEAD_BITS)-1:7*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_1[6*(2*BITS+OVERHEAD_BITS)-1:6*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_1[5*(2*BITS+OVERHEAD_BITS)-1:5*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_1[4*(2*BITS+OVERHEAD_BITS)-1:4*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_1[3*(2*BITS+OVERHEAD_BITS)-1:3*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_1[2*(2*BITS+OVERHEAD_BITS)-1:2*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_1[(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_1[(2*BITS+OVERHEAD_BITS)-1:(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsOddChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        otherWordsOddChannels_input_reg[12*BITS-1:0] <= {(12*BITS){1'b0}};
        write_address_otherWordsEvenChannels_reg <= first_row_writing_others + 6;
        case(results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= results_to_write_in_ram_2[18*(2*BITS+OVERHEAD_BITS)-1:18*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[30*BITS-1:29*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= results_to_write_in_ram_2[17*(2*BITS+OVERHEAD_BITS)-1:17*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[29*BITS-1:28*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= results_to_write_in_ram_2[16*(2*BITS+OVERHEAD_BITS)-1:16*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[28*BITS-1:27*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= results_to_write_in_ram_2[15*(2*BITS+OVERHEAD_BITS)-1:15*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[27*BITS-1:26*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= results_to_write_in_ram_2[14*(2*BITS+OVERHEAD_BITS)-1:14*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[26*BITS-1:25*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= results_to_write_in_ram_2[13*(2*BITS+OVERHEAD_BITS)-1:13*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[25*BITS-1:24*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= results_to_write_in_ram_2[12*(2*BITS+OVERHEAD_BITS)-1:12*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[24*BITS-1:23*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= results_to_write_in_ram_2[11*(2*BITS+OVERHEAD_BITS)-1:11*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[23*BITS-1:22*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= results_to_write_in_ram_2[10*(2*BITS+OVERHEAD_BITS)-1:10*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[22*BITS-1:21*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= results_to_write_in_ram_2[9*(2*BITS+OVERHEAD_BITS)-1:9*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[21*BITS-1:20*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= results_to_write_in_ram_2[8*(2*BITS+OVERHEAD_BITS)-1:8*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[20*BITS-1:19*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= results_to_write_in_ram_2[7*(2*BITS+OVERHEAD_BITS)-1:7*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[19*BITS-1:18*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= results_to_write_in_ram_2[6*(2*BITS+OVERHEAD_BITS)-1:6*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[18*BITS-1:17*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= results_to_write_in_ram_2[5*(2*BITS+OVERHEAD_BITS)-1:5*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[17*BITS-1:16*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= results_to_write_in_ram_2[4*(2*BITS+OVERHEAD_BITS)-1:4*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[16*BITS-1:15*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= results_to_write_in_ram_2[3*(2*BITS+OVERHEAD_BITS)-1:3*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[15*BITS-1:14*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= results_to_write_in_ram_2[2*(2*BITS+OVERHEAD_BITS)-1:2*(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[14*BITS-1:13*BITS] <= {BITS{1'b0}};
        endcase
        case(results_to_write_in_ram_2[(2*BITS+OVERHEAD_BITS)-1])
        0   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= results_to_write_in_ram_2[(2*BITS+OVERHEAD_BITS)-1:(2*BITS+OVERHEAD_BITS)-BITS];
        1   :   otherWordsEvenChannels_input_reg[13*BITS-1:12*BITS] <= {BITS{1'b0}};
        endcase
        otherWordsEvenChannels_input_reg[12*BITS-1:0] <= {(12*BITS){1'b0}};
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end    
  15 :  begin
        write_otherWordsOddChannels_reg <= 0;
        write_otherWordsEvenChannels_reg <= 0;
        first_row_writing_others <= first_row_writing_others + 49;
        counter_internal_phase_4 <= counter_internal_phase_4 + 1;
        end
  endcase
  
    if (start_to_output == 1)   
        begin
        case(counter_internal_phase_6)
        0   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[204*(2*BITS+OVERHEAD_BITS)-1:204*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[203*(2*BITS+OVERHEAD_BITS)-1:203*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[204*(2*BITS+OVERHEAD_BITS)-1:204*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[203*(2*BITS+OVERHEAD_BITS)-1:203*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase 
        1   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[202*(2*BITS+OVERHEAD_BITS)-1:202*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[201*(2*BITS+OVERHEAD_BITS)-1:201*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[202*(2*BITS+OVERHEAD_BITS)-1:202*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[201*(2*BITS+OVERHEAD_BITS)-1:201*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase       
        2   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[200*(2*BITS+OVERHEAD_BITS)-1:200*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[199*(2*BITS+OVERHEAD_BITS)-1:199*(2*BITS+OVERHEAD_BITS)-BITS]};  
                1    :   output_channels_reg <= {results_to_write_in_ram_2[200*(2*BITS+OVERHEAD_BITS)-1:200*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[199*(2*BITS+OVERHEAD_BITS)-1:199*(2*BITS+OVERHEAD_BITS)-BITS]};  
                endcase   
        3   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[198*(2*BITS+OVERHEAD_BITS)-1:198*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[197*(2*BITS+OVERHEAD_BITS)-1:197*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[198*(2*BITS+OVERHEAD_BITS)-1:198*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[197*(2*BITS+OVERHEAD_BITS)-1:197*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase   
        4   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[196*(2*BITS+OVERHEAD_BITS)-1:196*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[195*(2*BITS+OVERHEAD_BITS)-1:195*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[196*(2*BITS+OVERHEAD_BITS)-1:196*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[195*(2*BITS+OVERHEAD_BITS)-1:195*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase    
        5   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[194*(2*BITS+OVERHEAD_BITS)-1:194*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[193*(2*BITS+OVERHEAD_BITS)-1:193*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[194*(2*BITS+OVERHEAD_BITS)-1:194*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[193*(2*BITS+OVERHEAD_BITS)-1:193*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase 
        6   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[192*(2*BITS+OVERHEAD_BITS)-1:192*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[191*(2*BITS+OVERHEAD_BITS)-1:191*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[192*(2*BITS+OVERHEAD_BITS)-1:192*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[191*(2*BITS+OVERHEAD_BITS)-1:191*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase       
        7   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[190*(2*BITS+OVERHEAD_BITS)-1:190*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[189*(2*BITS+OVERHEAD_BITS)-1:189*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[190*(2*BITS+OVERHEAD_BITS)-1:190*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[189*(2*BITS+OVERHEAD_BITS)-1:189*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        8   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[188*(2*BITS+OVERHEAD_BITS)-1:188*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[187*(2*BITS+OVERHEAD_BITS)-1:187*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[188*(2*BITS+OVERHEAD_BITS)-1:188*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[187*(2*BITS+OVERHEAD_BITS)-1:187*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase   
        9   :   case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[186*(2*BITS+OVERHEAD_BITS)-1:186*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[185*(2*BITS+OVERHEAD_BITS)-1:185*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[186*(2*BITS+OVERHEAD_BITS)-1:186*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[185*(2*BITS+OVERHEAD_BITS)-1:185*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase  
        10   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[184*(2*BITS+OVERHEAD_BITS)-1:184*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[183*(2*BITS+OVERHEAD_BITS)-1:183*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[184*(2*BITS+OVERHEAD_BITS)-1:184*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[183*(2*BITS+OVERHEAD_BITS)-1:183*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase 
        11   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[182*(2*BITS+OVERHEAD_BITS)-1:182*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[181*(2*BITS+OVERHEAD_BITS)-1:181*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[182*(2*BITS+OVERHEAD_BITS)-1:182*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[181*(2*BITS+OVERHEAD_BITS)-1:181*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase       
        12   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[180*(2*BITS+OVERHEAD_BITS)-1:180*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[179*(2*BITS+OVERHEAD_BITS)-1:179*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[180*(2*BITS+OVERHEAD_BITS)-1:180*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[179*(2*BITS+OVERHEAD_BITS)-1:179*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase   
        13   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[178*(2*BITS+OVERHEAD_BITS)-1:178*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[177*(2*BITS+OVERHEAD_BITS)-1:177*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[178*(2*BITS+OVERHEAD_BITS)-1:178*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[177*(2*BITS+OVERHEAD_BITS)-1:177*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase   
        14   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[176*(2*BITS+OVERHEAD_BITS)-1:176*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[175*(2*BITS+OVERHEAD_BITS)-1:175*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[176*(2*BITS+OVERHEAD_BITS)-1:176*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[175*(2*BITS+OVERHEAD_BITS)-1:175*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase    
        15   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[174*(2*BITS+OVERHEAD_BITS)-1:174*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[173*(2*BITS+OVERHEAD_BITS)-1:173*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[174*(2*BITS+OVERHEAD_BITS)-1:174*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[173*(2*BITS+OVERHEAD_BITS)-1:173*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase 
        16   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[172*(2*BITS+OVERHEAD_BITS)-1:172*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[171*(2*BITS+OVERHEAD_BITS)-1:171*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[172*(2*BITS+OVERHEAD_BITS)-1:172*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[171*(2*BITS+OVERHEAD_BITS)-1:171*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase       
        17   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[170*(2*BITS+OVERHEAD_BITS)-1:170*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[169*(2*BITS+OVERHEAD_BITS)-1:169*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[170*(2*BITS+OVERHEAD_BITS)-1:170*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[169*(2*BITS+OVERHEAD_BITS)-1:169*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase   
        18   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[168*(2*BITS+OVERHEAD_BITS)-1:168*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[167*(2*BITS+OVERHEAD_BITS)-1:167*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[168*(2*BITS+OVERHEAD_BITS)-1:168*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[167*(2*BITS+OVERHEAD_BITS)-1:167*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        19   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[166*(2*BITS+OVERHEAD_BITS)-1:166*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[165*(2*BITS+OVERHEAD_BITS)-1:165*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[166*(2*BITS+OVERHEAD_BITS)-1:166*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[165*(2*BITS+OVERHEAD_BITS)-1:165*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase
        20   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[164*(2*BITS+OVERHEAD_BITS)-1:164*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[163*(2*BITS+OVERHEAD_BITS)-1:163*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[164*(2*BITS+OVERHEAD_BITS)-1:164*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[163*(2*BITS+OVERHEAD_BITS)-1:163*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase 
        21   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[162*(2*BITS+OVERHEAD_BITS)-1:162*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[161*(2*BITS+OVERHEAD_BITS)-1:161*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[162*(2*BITS+OVERHEAD_BITS)-1:162*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[161*(2*BITS+OVERHEAD_BITS)-1:161*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase       
        22   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[160*(2*BITS+OVERHEAD_BITS)-1:160*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[159*(2*BITS+OVERHEAD_BITS)-1:159*(2*BITS+OVERHEAD_BITS)-BITS]};  
                1    :   output_channels_reg <= {results_to_write_in_ram_2[160*(2*BITS+OVERHEAD_BITS)-1:160*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[159*(2*BITS+OVERHEAD_BITS)-1:159*(2*BITS+OVERHEAD_BITS)-BITS]};  
                endcase   
        23   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[158*(2*BITS+OVERHEAD_BITS)-1:158*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[157*(2*BITS+OVERHEAD_BITS)-1:157*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[158*(2*BITS+OVERHEAD_BITS)-1:158*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[157*(2*BITS+OVERHEAD_BITS)-1:157*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase   
        24   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[156*(2*BITS+OVERHEAD_BITS)-1:156*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[155*(2*BITS+OVERHEAD_BITS)-1:155*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[156*(2*BITS+OVERHEAD_BITS)-1:156*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[155*(2*BITS+OVERHEAD_BITS)-1:155*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase    
        25   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[154*(2*BITS+OVERHEAD_BITS)-1:154*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[153*(2*BITS+OVERHEAD_BITS)-1:153*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[154*(2*BITS+OVERHEAD_BITS)-1:154*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[153*(2*BITS+OVERHEAD_BITS)-1:153*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase 
        26   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[152*(2*BITS+OVERHEAD_BITS)-1:152*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[151*(2*BITS+OVERHEAD_BITS)-1:151*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[152*(2*BITS+OVERHEAD_BITS)-1:152*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[151*(2*BITS+OVERHEAD_BITS)-1:151*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase       
        27   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[150*(2*BITS+OVERHEAD_BITS)-1:150*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[149*(2*BITS+OVERHEAD_BITS)-1:149*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[150*(2*BITS+OVERHEAD_BITS)-1:150*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[149*(2*BITS+OVERHEAD_BITS)-1:149*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        28   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[148*(2*BITS+OVERHEAD_BITS)-1:148*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[147*(2*BITS+OVERHEAD_BITS)-1:147*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[148*(2*BITS+OVERHEAD_BITS)-1:148*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[147*(2*BITS+OVERHEAD_BITS)-1:147*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase  
        29   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[146*(2*BITS+OVERHEAD_BITS)-1:146*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[145*(2*BITS+OVERHEAD_BITS)-1:145*(2*BITS+OVERHEAD_BITS)-BITS]};  
                1    :   output_channels_reg <= {results_to_write_in_ram_2[146*(2*BITS+OVERHEAD_BITS)-1:146*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[145*(2*BITS+OVERHEAD_BITS)-1:145*(2*BITS+OVERHEAD_BITS)-BITS]};  
                endcase  
        30   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[144*(2*BITS+OVERHEAD_BITS)-1:144*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[143*(2*BITS+OVERHEAD_BITS)-1:143*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[144*(2*BITS+OVERHEAD_BITS)-1:144*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[143*(2*BITS+OVERHEAD_BITS)-1:143*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase 
        31   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[142*(2*BITS+OVERHEAD_BITS)-1:142*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[141*(2*BITS+OVERHEAD_BITS)-1:141*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[142*(2*BITS+OVERHEAD_BITS)-1:142*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[141*(2*BITS+OVERHEAD_BITS)-1:141*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase       
        32   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[140*(2*BITS+OVERHEAD_BITS)-1:140*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[139*(2*BITS+OVERHEAD_BITS)-1:139*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[140*(2*BITS+OVERHEAD_BITS)-1:140*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[139*(2*BITS+OVERHEAD_BITS)-1:139*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase   
        33   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[138*(2*BITS+OVERHEAD_BITS)-1:138*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[137*(2*BITS+OVERHEAD_BITS)-1:137*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[138*(2*BITS+OVERHEAD_BITS)-1:138*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[137*(2*BITS+OVERHEAD_BITS)-1:137*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase  
        34   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[136*(2*BITS+OVERHEAD_BITS)-1:136*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[135*(2*BITS+OVERHEAD_BITS)-1:135*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[136*(2*BITS+OVERHEAD_BITS)-1:136*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[135*(2*BITS+OVERHEAD_BITS)-1:135*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase    
        35   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[134*(2*BITS+OVERHEAD_BITS)-1:134*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[133*(2*BITS+OVERHEAD_BITS)-1:133*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[134*(2*BITS+OVERHEAD_BITS)-1:134*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[133*(2*BITS+OVERHEAD_BITS)-1:133*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase 
        36   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[132*(2*BITS+OVERHEAD_BITS)-1:132*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[131*(2*BITS+OVERHEAD_BITS)-1:131*(2*BITS+OVERHEAD_BITS)-BITS]}; 
                1    :   output_channels_reg <= {results_to_write_in_ram_2[132*(2*BITS+OVERHEAD_BITS)-1:132*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[131*(2*BITS+OVERHEAD_BITS)-1:131*(2*BITS+OVERHEAD_BITS)-BITS]}; 
                endcase       
        37   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[130*(2*BITS+OVERHEAD_BITS)-1:130*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[129*(2*BITS+OVERHEAD_BITS)-1:129*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[130*(2*BITS+OVERHEAD_BITS)-1:130*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[129*(2*BITS+OVERHEAD_BITS)-1:129*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase   
        38   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[128*(2*BITS+OVERHEAD_BITS)-1:128*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[127*(2*BITS+OVERHEAD_BITS)-1:127*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[128*(2*BITS+OVERHEAD_BITS)-1:128*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[127*(2*BITS+OVERHEAD_BITS)-1:127*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase   
        39   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[126*(2*BITS+OVERHEAD_BITS)-1:126*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[125*(2*BITS+OVERHEAD_BITS)-1:125*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[126*(2*BITS+OVERHEAD_BITS)-1:126*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[125*(2*BITS+OVERHEAD_BITS)-1:125*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase  
        40   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[124*(2*BITS+OVERHEAD_BITS)-1:124*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[123*(2*BITS+OVERHEAD_BITS)-1:123*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[124*(2*BITS+OVERHEAD_BITS)-1:124*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[123*(2*BITS+OVERHEAD_BITS)-1:123*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase 
        41   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[122*(2*BITS+OVERHEAD_BITS)-1:122*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[121*(2*BITS+OVERHEAD_BITS)-1:121*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[122*(2*BITS+OVERHEAD_BITS)-1:122*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[121*(2*BITS+OVERHEAD_BITS)-1:121*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase       
        42   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[120*(2*BITS+OVERHEAD_BITS)-1:120*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[119*(2*BITS+OVERHEAD_BITS)-1:119*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[120*(2*BITS+OVERHEAD_BITS)-1:120*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[119*(2*BITS+OVERHEAD_BITS)-1:119*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase   
        43   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[118*(2*BITS+OVERHEAD_BITS)-1:118*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[117*(2*BITS+OVERHEAD_BITS)-1:117*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[118*(2*BITS+OVERHEAD_BITS)-1:118*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[117*(2*BITS+OVERHEAD_BITS)-1:117*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        44   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[116*(2*BITS+OVERHEAD_BITS)-1:116*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[115*(2*BITS+OVERHEAD_BITS)-1:115*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[116*(2*BITS+OVERHEAD_BITS)-1:116*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[115*(2*BITS+OVERHEAD_BITS)-1:115*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase    
        45   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[114*(2*BITS+OVERHEAD_BITS)-1:114*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[113*(2*BITS+OVERHEAD_BITS)-1:113*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[114*(2*BITS+OVERHEAD_BITS)-1:114*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[113*(2*BITS+OVERHEAD_BITS)-1:113*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase 
        46   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[112*(2*BITS+OVERHEAD_BITS)-1:112*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[111*(2*BITS+OVERHEAD_BITS)-1:111*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[112*(2*BITS+OVERHEAD_BITS)-1:112*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[111*(2*BITS+OVERHEAD_BITS)-1:111*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase       
        47   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[110*(2*BITS+OVERHEAD_BITS)-1:110*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[109*(2*BITS+OVERHEAD_BITS)-1:109*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[110*(2*BITS+OVERHEAD_BITS)-1:110*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[109*(2*BITS+OVERHEAD_BITS)-1:109*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        48   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[108*(2*BITS+OVERHEAD_BITS)-1:108*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[107*(2*BITS+OVERHEAD_BITS)-1:107*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[108*(2*BITS+OVERHEAD_BITS)-1:108*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[107*(2*BITS+OVERHEAD_BITS)-1:107*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase   
        49   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[106*(2*BITS+OVERHEAD_BITS)-1:106*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[105*(2*BITS+OVERHEAD_BITS)-1:105*(2*BITS+OVERHEAD_BITS)-BITS]}; 
                1    :   output_channels_reg <= {results_to_write_in_ram_2[106*(2*BITS+OVERHEAD_BITS)-1:106*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[105*(2*BITS+OVERHEAD_BITS)-1:105*(2*BITS+OVERHEAD_BITS)-BITS]}; 
                endcase
        50   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[104*(2*BITS+OVERHEAD_BITS)-1:104*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[103*(2*BITS+OVERHEAD_BITS)-1:103*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[104*(2*BITS+OVERHEAD_BITS)-1:104*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[103*(2*BITS+OVERHEAD_BITS)-1:103*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase 
        51   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[102*(2*BITS+OVERHEAD_BITS)-1:102*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[101*(2*BITS+OVERHEAD_BITS)-1:101*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[102*(2*BITS+OVERHEAD_BITS)-1:102*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[101*(2*BITS+OVERHEAD_BITS)-1:101*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase      
        52   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[100*(2*BITS+OVERHEAD_BITS)-1:100*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[99*(2*BITS+OVERHEAD_BITS)-1:99*(2*BITS+OVERHEAD_BITS)-BITS]};  
                1    :   output_channels_reg <= {results_to_write_in_ram_2[100*(2*BITS+OVERHEAD_BITS)-1:100*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[99*(2*BITS+OVERHEAD_BITS)-1:99*(2*BITS+OVERHEAD_BITS)-BITS]};  
                endcase   
        53   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[98*(2*BITS+OVERHEAD_BITS)-1:98*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[97*(2*BITS+OVERHEAD_BITS)-1:97*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[98*(2*BITS+OVERHEAD_BITS)-1:98*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[97*(2*BITS+OVERHEAD_BITS)-1:97*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase   
        54   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[96*(2*BITS+OVERHEAD_BITS)-1:96*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[95*(2*BITS+OVERHEAD_BITS)-1:95*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[96*(2*BITS+OVERHEAD_BITS)-1:96*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[95*(2*BITS+OVERHEAD_BITS)-1:95*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase    
        55   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[94*(2*BITS+OVERHEAD_BITS)-1:94*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[93*(2*BITS+OVERHEAD_BITS)-1:93*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[94*(2*BITS+OVERHEAD_BITS)-1:94*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[93*(2*BITS+OVERHEAD_BITS)-1:93*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase 
        56   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[92*(2*BITS+OVERHEAD_BITS)-1:92*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[91*(2*BITS+OVERHEAD_BITS)-1:91*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[92*(2*BITS+OVERHEAD_BITS)-1:92*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[91*(2*BITS+OVERHEAD_BITS)-1:91*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase       
        57   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[90*(2*BITS+OVERHEAD_BITS)-1:90*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[89*(2*BITS+OVERHEAD_BITS)-1:89*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[90*(2*BITS+OVERHEAD_BITS)-1:90*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[89*(2*BITS+OVERHEAD_BITS)-1:89*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        58   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[88*(2*BITS+OVERHEAD_BITS)-1:88*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[87*(2*BITS+OVERHEAD_BITS)-1:87*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[88*(2*BITS+OVERHEAD_BITS)-1:88*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[87*(2*BITS+OVERHEAD_BITS)-1:87*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        59   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[86*(2*BITS+OVERHEAD_BITS)-1:86*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[85*(2*BITS+OVERHEAD_BITS)-1:85*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[86*(2*BITS+OVERHEAD_BITS)-1:86*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[85*(2*BITS+OVERHEAD_BITS)-1:85*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase
        60   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[84*(2*BITS+OVERHEAD_BITS)-1:84*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[83*(2*BITS+OVERHEAD_BITS)-1:83*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[84*(2*BITS+OVERHEAD_BITS)-1:84*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[83*(2*BITS+OVERHEAD_BITS)-1:83*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase 
        61   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[82*(2*BITS+OVERHEAD_BITS)-1:82*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[81*(2*BITS+OVERHEAD_BITS)-1:81*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[82*(2*BITS+OVERHEAD_BITS)-1:82*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[81*(2*BITS+OVERHEAD_BITS)-1:81*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase       
        62   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[80*(2*BITS+OVERHEAD_BITS)-1:80*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[79*(2*BITS+OVERHEAD_BITS)-1:79*(2*BITS+OVERHEAD_BITS)-BITS]};  
                1    :   output_channels_reg <= {results_to_write_in_ram_2[80*(2*BITS+OVERHEAD_BITS)-1:80*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[79*(2*BITS+OVERHEAD_BITS)-1:79*(2*BITS+OVERHEAD_BITS)-BITS]};  
                endcase   
        63   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[78*(2*BITS+OVERHEAD_BITS)-1:78*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[77*(2*BITS+OVERHEAD_BITS)-1:77*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[78*(2*BITS+OVERHEAD_BITS)-1:78*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[77*(2*BITS+OVERHEAD_BITS)-1:77*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        64   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[76*(2*BITS+OVERHEAD_BITS)-1:76*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[75*(2*BITS+OVERHEAD_BITS)-1:75*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[76*(2*BITS+OVERHEAD_BITS)-1:76*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[75*(2*BITS+OVERHEAD_BITS)-1:75*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase    
        65   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[74*(2*BITS+OVERHEAD_BITS)-1:74*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[73*(2*BITS+OVERHEAD_BITS)-1:73*(2*BITS+OVERHEAD_BITS)-BITS]};  
                1    :   output_channels_reg <= {results_to_write_in_ram_2[74*(2*BITS+OVERHEAD_BITS)-1:74*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[73*(2*BITS+OVERHEAD_BITS)-1:73*(2*BITS+OVERHEAD_BITS)-BITS]};  
                endcase 
        66   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[72*(2*BITS+OVERHEAD_BITS)-1:72*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[71*(2*BITS+OVERHEAD_BITS)-1:71*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[72*(2*BITS+OVERHEAD_BITS)-1:72*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[71*(2*BITS+OVERHEAD_BITS)-1:71*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase       
        67   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[70*(2*BITS+OVERHEAD_BITS)-1:70*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[69*(2*BITS+OVERHEAD_BITS)-1:69*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[70*(2*BITS+OVERHEAD_BITS)-1:70*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[69*(2*BITS+OVERHEAD_BITS)-1:69*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase   
        68   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[68*(2*BITS+OVERHEAD_BITS)-1:68*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[67*(2*BITS+OVERHEAD_BITS)-1:67*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[68*(2*BITS+OVERHEAD_BITS)-1:68*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[67*(2*BITS+OVERHEAD_BITS)-1:67*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase   
        69   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[66*(2*BITS+OVERHEAD_BITS)-1:66*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[65*(2*BITS+OVERHEAD_BITS)-1:65*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[66*(2*BITS+OVERHEAD_BITS)-1:66*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[65*(2*BITS+OVERHEAD_BITS)-1:65*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase
        70   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[64*(2*BITS+OVERHEAD_BITS)-1:64*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[63*(2*BITS+OVERHEAD_BITS)-1:63*(2*BITS+OVERHEAD_BITS)-BITS]}; 
                1    :   output_channels_reg <= {results_to_write_in_ram_2[64*(2*BITS+OVERHEAD_BITS)-1:64*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[63*(2*BITS+OVERHEAD_BITS)-1:63*(2*BITS+OVERHEAD_BITS)-BITS]}; 
                endcase 
        71   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[62*(2*BITS+OVERHEAD_BITS)-1:62*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[61*(2*BITS+OVERHEAD_BITS)-1:61*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[62*(2*BITS+OVERHEAD_BITS)-1:62*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[61*(2*BITS+OVERHEAD_BITS)-1:61*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase       
        72   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[60*(2*BITS+OVERHEAD_BITS)-1:60*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[59*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[60*(2*BITS+OVERHEAD_BITS)-1:60*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[59*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase   
        73   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[58*(2*BITS+OVERHEAD_BITS)-1:58*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[57*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[58*(2*BITS+OVERHEAD_BITS)-1:58*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[57*(2*BITS+OVERHEAD_BITS)-1:57*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        74   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[56*(2*BITS+OVERHEAD_BITS)-1:56*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[55*(2*BITS+OVERHEAD_BITS)-1:55*(2*BITS+OVERHEAD_BITS)-BITS]};  
                1    :   output_channels_reg <= {results_to_write_in_ram_2[56*(2*BITS+OVERHEAD_BITS)-1:56*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[55*(2*BITS+OVERHEAD_BITS)-1:55*(2*BITS+OVERHEAD_BITS)-BITS]};  
                endcase    
        75   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[54*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[53*(2*BITS+OVERHEAD_BITS)-1:53*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[54*(2*BITS+OVERHEAD_BITS)-1:54*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[53*(2*BITS+OVERHEAD_BITS)-1:53*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase 
        76   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[52*(2*BITS+OVERHEAD_BITS)-1:52*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[51*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[52*(2*BITS+OVERHEAD_BITS)-1:52*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[51*(2*BITS+OVERHEAD_BITS)-1:51*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase       
        77   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[50*(2*BITS+OVERHEAD_BITS)-1:50*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[49*(2*BITS+OVERHEAD_BITS)-1:49*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[50*(2*BITS+OVERHEAD_BITS)-1:50*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[49*(2*BITS+OVERHEAD_BITS)-1:49*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        78   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[48*(2*BITS+OVERHEAD_BITS)-1:48*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[47*(2*BITS+OVERHEAD_BITS)-1:47*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[48*(2*BITS+OVERHEAD_BITS)-1:48*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[47*(2*BITS+OVERHEAD_BITS)-1:47*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase   
        79   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[46*(2*BITS+OVERHEAD_BITS)-1:46*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[45*(2*BITS+OVERHEAD_BITS)-1:45*(2*BITS+OVERHEAD_BITS)-BITS]}; 
                1    :   output_channels_reg <= {results_to_write_in_ram_2[46*(2*BITS+OVERHEAD_BITS)-1:46*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[45*(2*BITS+OVERHEAD_BITS)-1:45*(2*BITS+OVERHEAD_BITS)-BITS]}; 
                endcase
        80   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[44*(2*BITS+OVERHEAD_BITS)-1:44*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[43*(2*BITS+OVERHEAD_BITS)-1:43*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[44*(2*BITS+OVERHEAD_BITS)-1:44*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[43*(2*BITS+OVERHEAD_BITS)-1:43*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase 
        81   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[42*(2*BITS+OVERHEAD_BITS)-1:42*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[41*(2*BITS+OVERHEAD_BITS)-1:41*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[42*(2*BITS+OVERHEAD_BITS)-1:42*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[41*(2*BITS+OVERHEAD_BITS)-1:41*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase       
        82   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[40*(2*BITS+OVERHEAD_BITS)-1:40*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[39*(2*BITS+OVERHEAD_BITS)-1:39*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[40*(2*BITS+OVERHEAD_BITS)-1:40*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[39*(2*BITS+OVERHEAD_BITS)-1:39*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase   
        83   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[38*(2*BITS+OVERHEAD_BITS)-1:38*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[37*(2*BITS+OVERHEAD_BITS)-1:37*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[38*(2*BITS+OVERHEAD_BITS)-1:38*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[37*(2*BITS+OVERHEAD_BITS)-1:37*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        84   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[36*(2*BITS+OVERHEAD_BITS)-1:36*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[35*(2*BITS+OVERHEAD_BITS)-1:35*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[36*(2*BITS+OVERHEAD_BITS)-1:36*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[35*(2*BITS+OVERHEAD_BITS)-1:35*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase    
        85   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[34*(2*BITS+OVERHEAD_BITS)-1:34*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[33*(2*BITS+OVERHEAD_BITS)-1:33*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[34*(2*BITS+OVERHEAD_BITS)-1:34*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[33*(2*BITS+OVERHEAD_BITS)-1:33*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase 
        86   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[32*(2*BITS+OVERHEAD_BITS)-1:32*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[31*(2*BITS+OVERHEAD_BITS)-1:31*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[32*(2*BITS+OVERHEAD_BITS)-1:32*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[31*(2*BITS+OVERHEAD_BITS)-1:31*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase       
        87   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[30*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[29*(2*BITS+OVERHEAD_BITS)-1:29*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[30*(2*BITS+OVERHEAD_BITS)-1:30*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[29*(2*BITS+OVERHEAD_BITS)-1:29*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        88   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[28*(2*BITS+OVERHEAD_BITS)-1:28*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[27*(2*BITS+OVERHEAD_BITS)-1:27*(2*BITS+OVERHEAD_BITS)-BITS]};      
                1    :   output_channels_reg <= {results_to_write_in_ram_2[28*(2*BITS+OVERHEAD_BITS)-1:28*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[27*(2*BITS+OVERHEAD_BITS)-1:27*(2*BITS+OVERHEAD_BITS)-BITS]};      
                endcase   
        89   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[26*(2*BITS+OVERHEAD_BITS)-1:26*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[25*(2*BITS+OVERHEAD_BITS)-1:25*(2*BITS+OVERHEAD_BITS)-BITS]};   
                1    :   output_channels_reg <= {results_to_write_in_ram_2[26*(2*BITS+OVERHEAD_BITS)-1:26*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[25*(2*BITS+OVERHEAD_BITS)-1:25*(2*BITS+OVERHEAD_BITS)-BITS]};   
                endcase
        90   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[24*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[23*(2*BITS+OVERHEAD_BITS)-1:23*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[24*(2*BITS+OVERHEAD_BITS)-1:24*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[23*(2*BITS+OVERHEAD_BITS)-1:23*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase 
        91   :  case(writing_row)                                                                     
                0    :   output_channels_reg <= {results_to_write_in_ram_1[22*(2*BITS+OVERHEAD_BITS)-1:22*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[21*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)-BITS]};    
                1    :   output_channels_reg <= {results_to_write_in_ram_2[22*(2*BITS+OVERHEAD_BITS)-1:22*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[21*(2*BITS+OVERHEAD_BITS)-1:21*(2*BITS+OVERHEAD_BITS)-BITS]};    
                endcase       
        92   :  case(writing_row)                                                                      
                0    :   output_channels_reg <= {results_to_write_in_ram_1[20*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_1[19*(2*BITS+OVERHEAD_BITS)-1:19*(2*BITS+OVERHEAD_BITS)-BITS]};     
                1    :   output_channels_reg <= {results_to_write_in_ram_2[20*(2*BITS+OVERHEAD_BITS)-1:20*(2*BITS+OVERHEAD_BITS)-BITS],results_to_write_in_ram_2[19*(2*BITS+OVERHEAD_BITS)-1:19*(2*BITS+OVERHEAD_BITS)-BITS]};     
                endcase   
        93   :  begin
                if (writing_row == 0)
                    begin
                    writing_row <= 1;
                    counter_internal_phase_6 <= 0;
                    end
                else
                    begin
                    counter_internal_phase_4 <= 16;
                    start_to_output <= 0;
                    end
                end
        endcase    
    end
    if (counter_internal_phase_6 < 93)
        begin
            counter_internal_phase_6 <= counter_internal_phase_6 + 1;
        end
    if (start_read_new_row == 1) 
        begin
            start_read_new_row <= 0; // te herschrijven bij integreren.
        end
    end
endmodule  
    
//if (start_read_new_row == 1'b1) 
//// Herschrijven, rekening houden met eerste klokcycli waar input binnenkomt. Dit test ik tijdens het integreren.
//    begin
//        start_read_new_row <= 1'b0;
//    end
//    
//if (start_to_output == 1)   
//    begin
//    case(counter_internal_phase_6)
//    9'b000000000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[192*BITS-1:190*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[192*BITS-1:190*BITS];
//                        endcase
//    9'b000000001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[190*BITS-1:188*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[190*BITS-1:188*BITS];
//                        endcase
//    9'b000000010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[188*BITS-1:186*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[188*BITS-1:186*BITS];
//                        endcase
//    9'b000000011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[186*BITS-1:184*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[186*BITS-1:184*BITS];
//                        endcase
//    9'b000000100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[184*BITS-1:182*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[184*BITS-1:182*BITS];
//                        endcase
//    9'b000000101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[182*BITS-1:180*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[182*BITS-1:180*BITS];
//                        endcase
//    9'b000000110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[180*BITS-1:178*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[180*BITS-1:178*BITS];
//                        endcase
//    9'b000000111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[178*BITS-1:176*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[178*BITS-1:176*BITS];
//                        endcase
//    9'b000001000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[176*BITS-1:174*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[176*BITS-1:174*BITS];
//                        endcase
//    9'b000001001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[174*BITS-1:172*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[174*BITS-1:172*BITS];
//                        endcase
//    9'b000001010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[172*BITS-1:170*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[172*BITS-1:170*BITS];
//                        endcase
//    9'b000001011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[170*BITS-1:168*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[170*BITS-1:168*BITS];
//                        endcase
//    9'b000001100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[168*BITS-1:166*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[168*BITS-1:166*BITS];
//                        endcase
//    9'b000001101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[166*BITS-1:164*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[166*BITS-1:164*BITS];
//                        endcase
//    9'b000001110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[164*BITS-1:162*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[164*BITS-1:162*BITS];
//                        endcase
//    9'b000001111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[162*BITS-1:160*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[162*BITS-1:160*BITS];
//                        endcase
//    9'b000010000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[160*BITS-1:158*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[160*BITS-1:158*BITS];
//                        endcase
//    9'b000010001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[158*BITS-1:156*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[158*BITS-1:156*BITS];
//                        endcase
//    9'b000010010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[156*BITS-1:154*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[156*BITS-1:154*BITS];
//                        endcase
//    9'b000010011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[154*BITS-1:152*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[154*BITS-1:152*BITS];
//                        endcase
//    9'b000010100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[152*BITS-1:150*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[152*BITS-1:150*BITS];
//                        endcase
//    9'b000010101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[150*BITS-1:148*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[150*BITS-1:148*BITS];
//                        endcase
//    9'b000010110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[148*BITS-1:146*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[148*BITS-1:146*BITS];
//                        endcase
//    9'b000010111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[146*BITS-1:144*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[146*BITS-1:144*BITS];
//                        endcase
//    9'b000011000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[144*BITS-1:142*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[144*BITS-1:142*BITS];
//                        endcase
//    9'b000011001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[142*BITS-1:140*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[142*BITS-1:140*BITS];
//                        endcase
//    9'b000011010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[140*BITS-1:138*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[140*BITS-1:138*BITS];
//                        endcase
//    9'b000011011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[138*BITS-1:136*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[138*BITS-1:136*BITS];
//                        endcase
//    9'b000011100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[136*BITS-1:134*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[136*BITS-1:134*BITS];
//                        endcase
//    9'b000011101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[134*BITS-1:132*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[134*BITS-1:132*BITS];
//                        endcase
//    9'b000011110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[132*BITS-1:130*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[132*BITS-1:130*BITS];
//                        endcase
//    9'b000011111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[130*BITS-1:128*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[130*BITS-1:128*BITS];
//                        endcase
//    9'b000100000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[128*BITS-1:126*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[128*BITS-1:126*BITS];
//                        endcase
//    9'b000100001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[126*BITS-1:124*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[126*BITS-1:124*BITS];
//                        endcase
//    9'b000100010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[124*BITS-1:122*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[124*BITS-1:122*BITS];
//                        endcase
//    9'b000100011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[122*BITS-1:120*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[122*BITS-1:120*BITS];
//                        endcase
//    9'b000100100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[120*BITS-1:118*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[120*BITS-1:118*BITS];
//                        endcase
//    9'b000100101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[118*BITS-1:116*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[118*BITS-1:116*BITS];
//                        endcase
//    9'b000100110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[116*BITS-1:114*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[116*BITS-1:114*BITS];
//                        endcase
//    9'b000100111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[114*BITS-1:112*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[114*BITS-1:112*BITS];
//                        endcase
//    9'b000101000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[112*BITS-1:110*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[112*BITS-1:110*BITS];
//                        endcase
//    9'b000101001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[110*BITS-1:108*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[110*BITS-1:108*BITS];
//                        endcase
//    9'b000101010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[108*BITS-1:106*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[108*BITS-1:106*BITS];
//                        endcase
//    9'b000101011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[106*BITS-1:104*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[106*BITS-1:104*BITS];
//                        endcase
//    9'b000101100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[104*BITS-1:102*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[104*BITS-1:102*BITS];
//                        endcase
//    9'b000101101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[102*BITS-1:100*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[102*BITS-1:100*BITS];
//                        endcase
//    9'b000101110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[100*BITS-1:98*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[100*BITS-1:98*BITS];
//                        endcase
//    9'b000101111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[98*BITS-1:96*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[98*BITS-1:96*BITS];
//                        endcase
//    9'b000110000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[96*BITS-1:94*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[96*BITS-1:94*BITS];
//                        endcase
//    9'b000110001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[94*BITS-1:92*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[94*BITS-1:92*BITS];
//                        endcase
//    9'b000110010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[92*BITS-1:90*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[92*BITS-1:90*BITS];
//                        endcase
//    9'b000110011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[90*BITS-1:88*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[90*BITS-1:88*BITS];
//                        endcase
//    9'b000110100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[88*BITS-1:86*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[88*BITS-1:86*BITS];
//                        endcase
//    9'b000110101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[86*BITS-1:84*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[86*BITS-1:84*BITS];
//                        endcase
//    9'b000110110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[84*BITS-1:82*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[84*BITS-1:82*BITS];
//                        endcase
//    9'b000110111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[82*BITS-1:80*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[82*BITS-1:80*BITS];
//                        endcase
//    9'b000111000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[80*BITS-1:78*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[80*BITS-1:78*BITS];
//                        endcase
//    9'b000111001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[78*BITS-1:76*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[78*BITS-1:76*BITS];
//                        endcase
//    9'b000111010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[76*BITS-1:74*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[76*BITS-1:74*BITS];
//                        endcase
//    9'b000111011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[74*BITS-1:72*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[74*BITS-1:72*BITS];
//                        endcase
//    9'b000111100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[72*BITS-1:70*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[72*BITS-1:70*BITS];
//                        endcase
//    9'b000111101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[70*BITS-1:68*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[70*BITS-1:68*BITS];
//                        endcase
//    9'b000111110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[68*BITS-1:66*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[68*BITS-1:66*BITS];
//                        endcase
//    9'b000111111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[66*BITS-1:64*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[66*BITS-1:64*BITS];
//                        endcase
//    9'b001000000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[64*BITS-1:62*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[64*BITS-1:62*BITS];
//                        endcase
//    9'b001000001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[62*BITS-1:60*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[62*BITS-1:60*BITS];
//                        endcase
//    9'b001000010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[60*BITS-1:58*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[60*BITS-1:58*BITS];
//                        endcase
//    9'b001000011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[58*BITS-1:56*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[58*BITS-1:56*BITS];
//                        endcase
//    9'b001000100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[56*BITS-1:54*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[56*BITS-1:54*BITS];
//                        endcase
//    9'b001000101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[54*BITS-1:52*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[54*BITS-1:52*BITS];
//                        endcase
//    9'b001000110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[52*BITS-1:50*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[52*BITS-1:50*BITS];
//                        endcase
//    9'b001000111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[50*BITS-1:48*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[50*BITS-1:48*BITS];
//                        endcase
//    9'b001001000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[48*BITS-1:46*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[48*BITS-1:46*BITS];
//                        endcase
//    9'b001001001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[46*BITS-1:44*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[46*BITS-1:44*BITS];
//                        endcase
//    9'b001001010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[44*BITS-1:42*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[44*BITS-1:42*BITS];
//                        endcase
//    9'b001001011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[42*BITS-1:40*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[42*BITS-1:40*BITS];
//                        endcase
//    9'b001001100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[40*BITS-1:38*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[40*BITS-1:38*BITS];
//                        endcase
//    9'b001001101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[38*BITS-1:36*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[38*BITS-1:36*BITS];
//                        endcase
//    9'b001001110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[36*BITS-1:34*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[36*BITS-1:34*BITS];
//                        endcase
//    9'b001001111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[34*BITS-1:32*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[34*BITS-1:32*BITS];
//                        endcase
//    9'b001010000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[32*BITS-1:30*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[32*BITS-1:30*BITS];
//                        endcase
//    9'b001010001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[30*BITS-1:28*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[30*BITS-1:28*BITS];
//                        endcase
//    9'b001010010    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[28*BITS-1:26*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[28*BITS-1:26*BITS];
//                        endcase
//    9'b001010011    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[26*BITS-1:24*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[26*BITS-1:24*BITS];
//                        endcase
//    9'b001010100    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[24*BITS-1:22*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[24*BITS-1:22*BITS];
//                        endcase
//    9'b001010101    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[22*BITS-1:20*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[22*BITS-1:20*BITS];
//                        endcase
//    9'b001010110    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[20*BITS-1:18*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[20*BITS-1:18*BITS];
//                        endcase
//    9'b001010111    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[18*BITS-1:16*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[18*BITS-1:16*BITS];
//                        endcase
//    9'b001011000    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[16*BITS-1:14*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[16*BITS-1:14*BITS];
//                        endcase
//    9'b001011001    :   case(writing_row)
//                        1'b0    :   output_channels_reg <= results_to_write_in_ram_1[14*BITS-1:12*BITS];
//                        1'b1    :   output_channels_reg <= results_to_write_in_ram_2[14*BITS-1:12*BITS];
//                        endcase
//    9'b001011010    :   begin
//                        if (writing_row == 0)
//                            begin
//                            writing_row <= 1;
//                            counter_internal_phase_6 <= 0;
//                            end
//                        else
//                            begin
//                            counter_internal_phase_4 <= 5'b11111;
//                            start_to_output <= 0;
//                            end
//                        end
//    endcase    
//    if (counter_internal_phase_6 < 90)
//        begin
//            counter_internal_phase_6 <= counter_internal_phase_6 + 1;
//        end
//    end
//end



//assign features = 
//{temp_in_1[66*BITS-1-0:51*BITS],
//temp_in_1[66*BITS-BITS-1:66*BITS-(FEATURES-KERNEL+2)*BITS],
//temp_in_1[66*BITS-2*BITS-1:66*BITS-(FEATURES-KERNEL+3)*BITS],
//temp_in_1[66*BITS-3*BITS-1:66*BITS-(FEATURES-KERNEL+4)*BITS],
//temp_in_1[66*BITS-4*BITS-1:66*BITS-(FEATURES-KERNEL+5)*BITS],
//temp_in_1[66*BITS-5*BITS-1:66*BITS-(FEATURES-KERNEL+6)*BITS],
//temp_in_1[66*BITS-6*BITS-1:66*BITS-(FEATURES-KERNEL+7)*BITS],
//temp_in_2[66*BITS-1:66*BITS-(FEATURES-KERNEL+1)*BITS],
//temp_in_2[66*BITS-BITS-1:66*BITS-(FEATURES-KERNEL+2)*BITS],
//temp_in_2[66*BITS-2*BITS-1:66*BITS-(FEATURES-KERNEL+3)*BITS],
//temp_in_2[66*BITS-3*BITS-1:66*BITS-(FEATURES-KERNEL+4)*BITS],
//temp_in_2[66*BITS-4*BITS-1:66*BITS-(FEATURES-KERNEL+5)*BITS],
//temp_in_2[66*BITS-5*BITS-1:66*BITS-(FEATURES-KERNEL+6)*BITS],
//temp_in_2[66*BITS-6*BITS-1:66*BITS-(FEATURES-KERNEL+7)*BITS],
//temp_in_1[66*BITS-15*BITS-1:66*BITS-(FEATURES-KERNEL+16)*BITS],
//temp_in_1[66*BITS-16*BITS-1:66*BITS-(FEATURES-KERNEL+17)*BITS],
//temp_in_1[66*BITS-17*BITS-1:66*BITS-(FEATURES-KERNEL+18)*BITS],
//temp_in_1[66*BITS-18*BITS-1:66*BITS-(FEATURES-KERNEL+19)*BITS],
//temp_in_1[66*BITS-19*BITS-1:66*BITS-(FEATURES-KERNEL+20)*BITS],
//temp_in_1[66*BITS-20*BITS-1:66*BITS-(FEATURES-KERNEL+21)*BITS],
//temp_in_1[66*BITS-21*BITS-1:66*BITS-(FEATURES-KERNEL+22)*BITS],
//temp_in_2[66*BITS-15*BITS-1:66*BITS-(FEATURES-KERNEL+16)*BITS],
//temp_in_2[66*BITS-16*BITS-1:66*BITS-(FEATURES-KERNEL+17)*BITS],
//temp_in_2[66*BITS-17*BITS-1:66*BITS-(FEATURES-KERNEL+18)*BITS],
//temp_in_2[66*BITS-18*BITS-1:66*BITS-(FEATURES-KERNEL+19)*BITS],
//temp_in_2[66*BITS-19*BITS-1:66*BITS-(FEATURES-KERNEL+20)*BITS],
//temp_in_2[66*BITS-20*BITS-1:66*BITS-(FEATURES-KERNEL+21)*BITS],
//temp_in_2[66*BITS-21*BITS-1:66*BITS-(FEATURES-KERNEL+22)*BITS],
//temp_in_1[66*BITS-1:66*BITS-(FEATURES-KERNEL+1)*BITS],
//temp_in_1[66*BITS-BITS-1:66*BITS-(FEATURES-KERNEL+2)*BITS],
//temp_in_1[66*BITS-2*BITS-1:66*BITS-(FEATURES-KERNEL+3)*BITS],
//temp_in_1[66*BITS-3*BITS-1:66*BITS-(FEATURES-KERNEL+4)*BITS],
//temp_in_1[66*BITS-4*BITS-1:66*BITS-(FEATURES-KERNEL+5)*BITS],
//temp_in_1[66*BITS-5*BITS-1:66*BITS-(FEATURES-KERNEL+6)*BITS],
//temp_in_1[66*BITS-6*BITS-1:66*BITS-(FEATURES-KERNEL+7)*BITS],
//temp_in_2[66*BITS-1:66*BITS-(FEATURES-KERNEL+1)*BITS],
//temp_in_2[66*BITS-BITS-1:66*BITS-(FEATURES-KERNEL+2)*BITS],
//temp_in_2[66*BITS-2*BITS-1:66*BITS-(FEATURES-KERNEL+3)*BITS],
//temp_in_2[66*BITS-3*BITS-1:66*BITS-(FEATURES-KERNEL+4)*BITS],
//temp_in_2[66*BITS-4*BITS-1:66*BITS-(FEATURES-KERNEL+5)*BITS],
//temp_in_2[66*BITS-5*BITS-1:66*BITS-(FEATURES-KERNEL+6)*BITS],
//temp_in_2[66*BITS-6*BITS-1:66*BITS-(FEATURES-KERNEL+7)*BITS],
//temp_in_1[66*BITS-15*BITS-1:66*BITS-(FEATURES-KERNEL+16)*BITS],
//temp_in_1[66*BITS-16*BITS-1:66*BITS-(FEATURES-KERNEL+17)*BITS],
//temp_in_1[66*BITS-17*BITS-1:66*BITS-(FEATURES-KERNEL+18)*BITS],
//temp_in_1[66*BITS-18*BITS-1:66*BITS-(FEATURES-KERNEL+19)*BITS],
//temp_in_1[66*BITS-19*BITS-1:66*BITS-(FEATURES-KERNEL+20)*BITS],
//temp_in_1[66*BITS-20*BITS-1:66*BITS-(FEATURES-KERNEL+21)*BITS],
//temp_in_1[66*BITS-21*BITS-1:66*BITS-(FEATURES-KERNEL+22)*BITS],
//temp_in_2[66*BITS-15*BITS-1:66*BITS-(FEATURES-KERNEL+16)*BITS],
//temp_in_2[66*BITS-16*BITS-1:66*BITS-(FEATURES-KERNEL+17)*BITS],
//temp_in_2[66*BITS-17*BITS-1:66*BITS-(FEATURES-KERNEL+18)*BITS],
//temp_in_2[66*BITS-18*BITS-1:66*BITS-(FEATURES-KERNEL+19)*BITS],
//temp_in_2[66*BITS-19*BITS-1:66*BITS-(FEATURES-KERNEL+20)*BITS],
//temp_in_2[66*BITS-20*BITS-1:66*BITS-(FEATURES-KERNEL+21)*BITS],
//temp_in_2[66*BITS-21*BITS-1:66*BITS-(FEATURES-KERNEL+22)*BITS]
//    };

  

